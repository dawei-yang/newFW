-- ***** IRSX_store_cell model *****
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY T7_store_cell IS
PORT
(
   nramp : IN std_logic;
   STR : IN std_logic;
   PIXin : IN std_logic_vector(11 downto 0);
   SHout : OUT std_logic := 'Z'
);
END T7_store_cell;

ARCHITECTURE behavioral of T7_store_cell is
SIGNAL StoredData : std_logic_vector(11 downto 0);
SIGNAL Z : std_logic;
begin
process(PIXin, nramp, STR, Z)
--adjust these according to gcc_clk and related stuff
constant delay1 : time := 4 ns; -- depends on delays in gcc
constant delay_incr : time := 8 ns; -- half of gcc period
begin
if STR = '1' then StoredData <= PIXin;
end if;
-- SHout needs to go low, then high, otherwise dff doesn't work
-- Z used to reset everything after all digitizing done, not sure if necessary
if Z = '1' then 
	SHout <= 'Z';
	Z <= '0' after delay_incr;
end if;
if falling_edge(nramp) then 
	SHout <= '0';
	Z <= '1' after delay1 + 4096*delay_incr;
end if;

if nramp = '0' and StoredData = "000000000000" then SHout <= '1' after delay1;
elsif nramp = '0' and StoredData = "000000000001" then SHout <= '1' after delay1 + 1*delay_incr;
elsif nramp = '0' and StoredData = "000000000010" then SHout <= '1' after delay1 + 2*delay_incr;
elsif nramp = '0' and StoredData = "000000000011" then SHout <= '1' after delay1 + 3*delay_incr;
elsif nramp = '0' and StoredData = "000000000100" then SHout <= '1' after delay1 + 4*delay_incr;
elsif nramp = '0' and StoredData = "000000000101" then SHout <= '1' after delay1 + 5*delay_incr;
elsif nramp = '0' and StoredData = "000000000110" then SHout <= '1' after delay1 + 6*delay_incr;
elsif nramp = '0' and StoredData = "000000000111" then SHout <= '1' after delay1 + 7*delay_incr;
elsif nramp = '0' and StoredData = "000000001000" then SHout <= '1' after delay1 + 8*delay_incr;
elsif nramp = '0' and StoredData = "000000001001" then SHout <= '1' after delay1 + 9*delay_incr;
elsif nramp = '0' and StoredData = "000000001010" then SHout <= '1' after delay1 + 10*delay_incr;
elsif nramp = '0' and StoredData = "000000001011" then SHout <= '1' after delay1 + 11*delay_incr;
elsif nramp = '0' and StoredData = "000000001100" then SHout <= '1' after delay1 + 12*delay_incr;
elsif nramp = '0' and StoredData = "000000001101" then SHout <= '1' after delay1 + 13*delay_incr;
elsif nramp = '0' and StoredData = "000000001110" then SHout <= '1' after delay1 + 14*delay_incr;
elsif nramp = '0' and StoredData = "000000001111" then SHout <= '1' after delay1 + 15*delay_incr;
elsif nramp = '0' and StoredData = "000000010000" then SHout <= '1' after delay1 + 16*delay_incr;
elsif nramp = '0' and StoredData = "000000010001" then SHout <= '1' after delay1 + 17*delay_incr;
elsif nramp = '0' and StoredData = "000000010010" then SHout <= '1' after delay1 + 18*delay_incr;
elsif nramp = '0' and StoredData = "000000010011" then SHout <= '1' after delay1 + 19*delay_incr;
elsif nramp = '0' and StoredData = "000000010100" then SHout <= '1' after delay1 + 20*delay_incr;
elsif nramp = '0' and StoredData = "000000010101" then SHout <= '1' after delay1 + 21*delay_incr;
elsif nramp = '0' and StoredData = "000000010110" then SHout <= '1' after delay1 + 22*delay_incr;
elsif nramp = '0' and StoredData = "000000010111" then SHout <= '1' after delay1 + 23*delay_incr;
elsif nramp = '0' and StoredData = "000000011000" then SHout <= '1' after delay1 + 24*delay_incr;
elsif nramp = '0' and StoredData = "000000011001" then SHout <= '1' after delay1 + 25*delay_incr;
elsif nramp = '0' and StoredData = "000000011010" then SHout <= '1' after delay1 + 26*delay_incr;
elsif nramp = '0' and StoredData = "000000011011" then SHout <= '1' after delay1 + 27*delay_incr;
elsif nramp = '0' and StoredData = "000000011100" then SHout <= '1' after delay1 + 28*delay_incr;
elsif nramp = '0' and StoredData = "000000011101" then SHout <= '1' after delay1 + 29*delay_incr;
elsif nramp = '0' and StoredData = "000000011110" then SHout <= '1' after delay1 + 30*delay_incr;
elsif nramp = '0' and StoredData = "000000011111" then SHout <= '1' after delay1 + 31*delay_incr;
elsif nramp = '0' and StoredData = "000000100000" then SHout <= '1' after delay1 + 32*delay_incr;
elsif nramp = '0' and StoredData = "000000100001" then SHout <= '1' after delay1 + 33*delay_incr;
elsif nramp = '0' and StoredData = "000000100010" then SHout <= '1' after delay1 + 34*delay_incr;
elsif nramp = '0' and StoredData = "000000100011" then SHout <= '1' after delay1 + 35*delay_incr;
elsif nramp = '0' and StoredData = "000000100100" then SHout <= '1' after delay1 + 36*delay_incr;
elsif nramp = '0' and StoredData = "000000100101" then SHout <= '1' after delay1 + 37*delay_incr;
elsif nramp = '0' and StoredData = "000000100110" then SHout <= '1' after delay1 + 38*delay_incr;
elsif nramp = '0' and StoredData = "000000100111" then SHout <= '1' after delay1 + 39*delay_incr;
elsif nramp = '0' and StoredData = "000000101000" then SHout <= '1' after delay1 + 40*delay_incr;
elsif nramp = '0' and StoredData = "000000101001" then SHout <= '1' after delay1 + 41*delay_incr;
elsif nramp = '0' and StoredData = "000000101010" then SHout <= '1' after delay1 + 42*delay_incr;
elsif nramp = '0' and StoredData = "000000101011" then SHout <= '1' after delay1 + 43*delay_incr;
elsif nramp = '0' and StoredData = "000000101100" then SHout <= '1' after delay1 + 44*delay_incr;
elsif nramp = '0' and StoredData = "000000101101" then SHout <= '1' after delay1 + 45*delay_incr;
elsif nramp = '0' and StoredData = "000000101110" then SHout <= '1' after delay1 + 46*delay_incr;
elsif nramp = '0' and StoredData = "000000101111" then SHout <= '1' after delay1 + 47*delay_incr;
elsif nramp = '0' and StoredData = "000000110000" then SHout <= '1' after delay1 + 48*delay_incr;
elsif nramp = '0' and StoredData = "000000110001" then SHout <= '1' after delay1 + 49*delay_incr;
elsif nramp = '0' and StoredData = "000000110010" then SHout <= '1' after delay1 + 50*delay_incr;
elsif nramp = '0' and StoredData = "000000110011" then SHout <= '1' after delay1 + 51*delay_incr;
elsif nramp = '0' and StoredData = "000000110100" then SHout <= '1' after delay1 + 52*delay_incr;
elsif nramp = '0' and StoredData = "000000110101" then SHout <= '1' after delay1 + 53*delay_incr;
elsif nramp = '0' and StoredData = "000000110110" then SHout <= '1' after delay1 + 54*delay_incr;
elsif nramp = '0' and StoredData = "000000110111" then SHout <= '1' after delay1 + 55*delay_incr;
elsif nramp = '0' and StoredData = "000000111000" then SHout <= '1' after delay1 + 56*delay_incr;
elsif nramp = '0' and StoredData = "000000111001" then SHout <= '1' after delay1 + 57*delay_incr;
elsif nramp = '0' and StoredData = "000000111010" then SHout <= '1' after delay1 + 58*delay_incr;
elsif nramp = '0' and StoredData = "000000111011" then SHout <= '1' after delay1 + 59*delay_incr;
elsif nramp = '0' and StoredData = "000000111100" then SHout <= '1' after delay1 + 60*delay_incr;
elsif nramp = '0' and StoredData = "000000111101" then SHout <= '1' after delay1 + 61*delay_incr;
elsif nramp = '0' and StoredData = "000000111110" then SHout <= '1' after delay1 + 62*delay_incr;
elsif nramp = '0' and StoredData = "000000111111" then SHout <= '1' after delay1 + 63*delay_incr;
elsif nramp = '0' and StoredData = "000001000000" then SHout <= '1' after delay1 + 64*delay_incr;
elsif nramp = '0' and StoredData = "000001000001" then SHout <= '1' after delay1 + 65*delay_incr;
elsif nramp = '0' and StoredData = "000001000010" then SHout <= '1' after delay1 + 66*delay_incr;
elsif nramp = '0' and StoredData = "000001000011" then SHout <= '1' after delay1 + 67*delay_incr;
elsif nramp = '0' and StoredData = "000001000100" then SHout <= '1' after delay1 + 68*delay_incr;
elsif nramp = '0' and StoredData = "000001000101" then SHout <= '1' after delay1 + 69*delay_incr;
elsif nramp = '0' and StoredData = "000001000110" then SHout <= '1' after delay1 + 70*delay_incr;
elsif nramp = '0' and StoredData = "000001000111" then SHout <= '1' after delay1 + 71*delay_incr;
elsif nramp = '0' and StoredData = "000001001000" then SHout <= '1' after delay1 + 72*delay_incr;
elsif nramp = '0' and StoredData = "000001001001" then SHout <= '1' after delay1 + 73*delay_incr;
elsif nramp = '0' and StoredData = "000001001010" then SHout <= '1' after delay1 + 74*delay_incr;
elsif nramp = '0' and StoredData = "000001001011" then SHout <= '1' after delay1 + 75*delay_incr;
elsif nramp = '0' and StoredData = "000001001100" then SHout <= '1' after delay1 + 76*delay_incr;
elsif nramp = '0' and StoredData = "000001001101" then SHout <= '1' after delay1 + 77*delay_incr;
elsif nramp = '0' and StoredData = "000001001110" then SHout <= '1' after delay1 + 78*delay_incr;
elsif nramp = '0' and StoredData = "000001001111" then SHout <= '1' after delay1 + 79*delay_incr;
elsif nramp = '0' and StoredData = "000001010000" then SHout <= '1' after delay1 + 80*delay_incr;
elsif nramp = '0' and StoredData = "000001010001" then SHout <= '1' after delay1 + 81*delay_incr;
elsif nramp = '0' and StoredData = "000001010010" then SHout <= '1' after delay1 + 82*delay_incr;
elsif nramp = '0' and StoredData = "000001010011" then SHout <= '1' after delay1 + 83*delay_incr;
elsif nramp = '0' and StoredData = "000001010100" then SHout <= '1' after delay1 + 84*delay_incr;
elsif nramp = '0' and StoredData = "000001010101" then SHout <= '1' after delay1 + 85*delay_incr;
elsif nramp = '0' and StoredData = "000001010110" then SHout <= '1' after delay1 + 86*delay_incr;
elsif nramp = '0' and StoredData = "000001010111" then SHout <= '1' after delay1 + 87*delay_incr;
elsif nramp = '0' and StoredData = "000001011000" then SHout <= '1' after delay1 + 88*delay_incr;
elsif nramp = '0' and StoredData = "000001011001" then SHout <= '1' after delay1 + 89*delay_incr;
elsif nramp = '0' and StoredData = "000001011010" then SHout <= '1' after delay1 + 90*delay_incr;
elsif nramp = '0' and StoredData = "000001011011" then SHout <= '1' after delay1 + 91*delay_incr;
elsif nramp = '0' and StoredData = "000001011100" then SHout <= '1' after delay1 + 92*delay_incr;
elsif nramp = '0' and StoredData = "000001011101" then SHout <= '1' after delay1 + 93*delay_incr;
elsif nramp = '0' and StoredData = "000001011110" then SHout <= '1' after delay1 + 94*delay_incr;
elsif nramp = '0' and StoredData = "000001011111" then SHout <= '1' after delay1 + 95*delay_incr;
elsif nramp = '0' and StoredData = "000001100000" then SHout <= '1' after delay1 + 96*delay_incr;
elsif nramp = '0' and StoredData = "000001100001" then SHout <= '1' after delay1 + 97*delay_incr;
elsif nramp = '0' and StoredData = "000001100010" then SHout <= '1' after delay1 + 98*delay_incr;
elsif nramp = '0' and StoredData = "000001100011" then SHout <= '1' after delay1 + 99*delay_incr;
elsif nramp = '0' and StoredData = "000001100100" then SHout <= '1' after delay1 + 100*delay_incr;
elsif nramp = '0' and StoredData = "000001100101" then SHout <= '1' after delay1 + 101*delay_incr;
elsif nramp = '0' and StoredData = "000001100110" then SHout <= '1' after delay1 + 102*delay_incr;
elsif nramp = '0' and StoredData = "000001100111" then SHout <= '1' after delay1 + 103*delay_incr;
elsif nramp = '0' and StoredData = "000001101000" then SHout <= '1' after delay1 + 104*delay_incr;
elsif nramp = '0' and StoredData = "000001101001" then SHout <= '1' after delay1 + 105*delay_incr;
elsif nramp = '0' and StoredData = "000001101010" then SHout <= '1' after delay1 + 106*delay_incr;
elsif nramp = '0' and StoredData = "000001101011" then SHout <= '1' after delay1 + 107*delay_incr;
elsif nramp = '0' and StoredData = "000001101100" then SHout <= '1' after delay1 + 108*delay_incr;
elsif nramp = '0' and StoredData = "000001101101" then SHout <= '1' after delay1 + 109*delay_incr;
elsif nramp = '0' and StoredData = "000001101110" then SHout <= '1' after delay1 + 110*delay_incr;
elsif nramp = '0' and StoredData = "000001101111" then SHout <= '1' after delay1 + 111*delay_incr;
elsif nramp = '0' and StoredData = "000001110000" then SHout <= '1' after delay1 + 112*delay_incr;
elsif nramp = '0' and StoredData = "000001110001" then SHout <= '1' after delay1 + 113*delay_incr;
elsif nramp = '0' and StoredData = "000001110010" then SHout <= '1' after delay1 + 114*delay_incr;
elsif nramp = '0' and StoredData = "000001110011" then SHout <= '1' after delay1 + 115*delay_incr;
elsif nramp = '0' and StoredData = "000001110100" then SHout <= '1' after delay1 + 116*delay_incr;
elsif nramp = '0' and StoredData = "000001110101" then SHout <= '1' after delay1 + 117*delay_incr;
elsif nramp = '0' and StoredData = "000001110110" then SHout <= '1' after delay1 + 118*delay_incr;
elsif nramp = '0' and StoredData = "000001110111" then SHout <= '1' after delay1 + 119*delay_incr;
elsif nramp = '0' and StoredData = "000001111000" then SHout <= '1' after delay1 + 120*delay_incr;
elsif nramp = '0' and StoredData = "000001111001" then SHout <= '1' after delay1 + 121*delay_incr;
elsif nramp = '0' and StoredData = "000001111010" then SHout <= '1' after delay1 + 122*delay_incr;
elsif nramp = '0' and StoredData = "000001111011" then SHout <= '1' after delay1 + 123*delay_incr;
elsif nramp = '0' and StoredData = "000001111100" then SHout <= '1' after delay1 + 124*delay_incr;
elsif nramp = '0' and StoredData = "000001111101" then SHout <= '1' after delay1 + 125*delay_incr;
elsif nramp = '0' and StoredData = "000001111110" then SHout <= '1' after delay1 + 126*delay_incr;
elsif nramp = '0' and StoredData = "000001111111" then SHout <= '1' after delay1 + 127*delay_incr;
elsif nramp = '0' and StoredData = "000010000000" then SHout <= '1' after delay1 + 128*delay_incr;
elsif nramp = '0' and StoredData = "000010000001" then SHout <= '1' after delay1 + 129*delay_incr;
elsif nramp = '0' and StoredData = "000010000010" then SHout <= '1' after delay1 + 130*delay_incr;
elsif nramp = '0' and StoredData = "000010000011" then SHout <= '1' after delay1 + 131*delay_incr;
elsif nramp = '0' and StoredData = "000010000100" then SHout <= '1' after delay1 + 132*delay_incr;
elsif nramp = '0' and StoredData = "000010000101" then SHout <= '1' after delay1 + 133*delay_incr;
elsif nramp = '0' and StoredData = "000010000110" then SHout <= '1' after delay1 + 134*delay_incr;
elsif nramp = '0' and StoredData = "000010000111" then SHout <= '1' after delay1 + 135*delay_incr;
elsif nramp = '0' and StoredData = "000010001000" then SHout <= '1' after delay1 + 136*delay_incr;
elsif nramp = '0' and StoredData = "000010001001" then SHout <= '1' after delay1 + 137*delay_incr;
elsif nramp = '0' and StoredData = "000010001010" then SHout <= '1' after delay1 + 138*delay_incr;
elsif nramp = '0' and StoredData = "000010001011" then SHout <= '1' after delay1 + 139*delay_incr;
elsif nramp = '0' and StoredData = "000010001100" then SHout <= '1' after delay1 + 140*delay_incr;
elsif nramp = '0' and StoredData = "000010001101" then SHout <= '1' after delay1 + 141*delay_incr;
elsif nramp = '0' and StoredData = "000010001110" then SHout <= '1' after delay1 + 142*delay_incr;
elsif nramp = '0' and StoredData = "000010001111" then SHout <= '1' after delay1 + 143*delay_incr;
elsif nramp = '0' and StoredData = "000010010000" then SHout <= '1' after delay1 + 144*delay_incr;
elsif nramp = '0' and StoredData = "000010010001" then SHout <= '1' after delay1 + 145*delay_incr;
elsif nramp = '0' and StoredData = "000010010010" then SHout <= '1' after delay1 + 146*delay_incr;
elsif nramp = '0' and StoredData = "000010010011" then SHout <= '1' after delay1 + 147*delay_incr;
elsif nramp = '0' and StoredData = "000010010100" then SHout <= '1' after delay1 + 148*delay_incr;
elsif nramp = '0' and StoredData = "000010010101" then SHout <= '1' after delay1 + 149*delay_incr;
elsif nramp = '0' and StoredData = "000010010110" then SHout <= '1' after delay1 + 150*delay_incr;
elsif nramp = '0' and StoredData = "000010010111" then SHout <= '1' after delay1 + 151*delay_incr;
elsif nramp = '0' and StoredData = "000010011000" then SHout <= '1' after delay1 + 152*delay_incr;
elsif nramp = '0' and StoredData = "000010011001" then SHout <= '1' after delay1 + 153*delay_incr;
elsif nramp = '0' and StoredData = "000010011010" then SHout <= '1' after delay1 + 154*delay_incr;
elsif nramp = '0' and StoredData = "000010011011" then SHout <= '1' after delay1 + 155*delay_incr;
elsif nramp = '0' and StoredData = "000010011100" then SHout <= '1' after delay1 + 156*delay_incr;
elsif nramp = '0' and StoredData = "000010011101" then SHout <= '1' after delay1 + 157*delay_incr;
elsif nramp = '0' and StoredData = "000010011110" then SHout <= '1' after delay1 + 158*delay_incr;
elsif nramp = '0' and StoredData = "000010011111" then SHout <= '1' after delay1 + 159*delay_incr;
elsif nramp = '0' and StoredData = "000010100000" then SHout <= '1' after delay1 + 160*delay_incr;
elsif nramp = '0' and StoredData = "000010100001" then SHout <= '1' after delay1 + 161*delay_incr;
elsif nramp = '0' and StoredData = "000010100010" then SHout <= '1' after delay1 + 162*delay_incr;
elsif nramp = '0' and StoredData = "000010100011" then SHout <= '1' after delay1 + 163*delay_incr;
elsif nramp = '0' and StoredData = "000010100100" then SHout <= '1' after delay1 + 164*delay_incr;
elsif nramp = '0' and StoredData = "000010100101" then SHout <= '1' after delay1 + 165*delay_incr;
elsif nramp = '0' and StoredData = "000010100110" then SHout <= '1' after delay1 + 166*delay_incr;
elsif nramp = '0' and StoredData = "000010100111" then SHout <= '1' after delay1 + 167*delay_incr;
elsif nramp = '0' and StoredData = "000010101000" then SHout <= '1' after delay1 + 168*delay_incr;
elsif nramp = '0' and StoredData = "000010101001" then SHout <= '1' after delay1 + 169*delay_incr;
elsif nramp = '0' and StoredData = "000010101010" then SHout <= '1' after delay1 + 170*delay_incr;
elsif nramp = '0' and StoredData = "000010101011" then SHout <= '1' after delay1 + 171*delay_incr;
elsif nramp = '0' and StoredData = "000010101100" then SHout <= '1' after delay1 + 172*delay_incr;
elsif nramp = '0' and StoredData = "000010101101" then SHout <= '1' after delay1 + 173*delay_incr;
elsif nramp = '0' and StoredData = "000010101110" then SHout <= '1' after delay1 + 174*delay_incr;
elsif nramp = '0' and StoredData = "000010101111" then SHout <= '1' after delay1 + 175*delay_incr;
elsif nramp = '0' and StoredData = "000010110000" then SHout <= '1' after delay1 + 176*delay_incr;
elsif nramp = '0' and StoredData = "000010110001" then SHout <= '1' after delay1 + 177*delay_incr;
elsif nramp = '0' and StoredData = "000010110010" then SHout <= '1' after delay1 + 178*delay_incr;
elsif nramp = '0' and StoredData = "000010110011" then SHout <= '1' after delay1 + 179*delay_incr;
elsif nramp = '0' and StoredData = "000010110100" then SHout <= '1' after delay1 + 180*delay_incr;
elsif nramp = '0' and StoredData = "000010110101" then SHout <= '1' after delay1 + 181*delay_incr;
elsif nramp = '0' and StoredData = "000010110110" then SHout <= '1' after delay1 + 182*delay_incr;
elsif nramp = '0' and StoredData = "000010110111" then SHout <= '1' after delay1 + 183*delay_incr;
elsif nramp = '0' and StoredData = "000010111000" then SHout <= '1' after delay1 + 184*delay_incr;
elsif nramp = '0' and StoredData = "000010111001" then SHout <= '1' after delay1 + 185*delay_incr;
elsif nramp = '0' and StoredData = "000010111010" then SHout <= '1' after delay1 + 186*delay_incr;
elsif nramp = '0' and StoredData = "000010111011" then SHout <= '1' after delay1 + 187*delay_incr;
elsif nramp = '0' and StoredData = "000010111100" then SHout <= '1' after delay1 + 188*delay_incr;
elsif nramp = '0' and StoredData = "000010111101" then SHout <= '1' after delay1 + 189*delay_incr;
elsif nramp = '0' and StoredData = "000010111110" then SHout <= '1' after delay1 + 190*delay_incr;
elsif nramp = '0' and StoredData = "000010111111" then SHout <= '1' after delay1 + 191*delay_incr;
elsif nramp = '0' and StoredData = "000011000000" then SHout <= '1' after delay1 + 192*delay_incr;
elsif nramp = '0' and StoredData = "000011000001" then SHout <= '1' after delay1 + 193*delay_incr;
elsif nramp = '0' and StoredData = "000011000010" then SHout <= '1' after delay1 + 194*delay_incr;
elsif nramp = '0' and StoredData = "000011000011" then SHout <= '1' after delay1 + 195*delay_incr;
elsif nramp = '0' and StoredData = "000011000100" then SHout <= '1' after delay1 + 196*delay_incr;
elsif nramp = '0' and StoredData = "000011000101" then SHout <= '1' after delay1 + 197*delay_incr;
elsif nramp = '0' and StoredData = "000011000110" then SHout <= '1' after delay1 + 198*delay_incr;
elsif nramp = '0' and StoredData = "000011000111" then SHout <= '1' after delay1 + 199*delay_incr;
elsif nramp = '0' and StoredData = "000011001000" then SHout <= '1' after delay1 + 200*delay_incr;
elsif nramp = '0' and StoredData = "000011001001" then SHout <= '1' after delay1 + 201*delay_incr;
elsif nramp = '0' and StoredData = "000011001010" then SHout <= '1' after delay1 + 202*delay_incr;
elsif nramp = '0' and StoredData = "000011001011" then SHout <= '1' after delay1 + 203*delay_incr;
elsif nramp = '0' and StoredData = "000011001100" then SHout <= '1' after delay1 + 204*delay_incr;
elsif nramp = '0' and StoredData = "000011001101" then SHout <= '1' after delay1 + 205*delay_incr;
elsif nramp = '0' and StoredData = "000011001110" then SHout <= '1' after delay1 + 206*delay_incr;
elsif nramp = '0' and StoredData = "000011001111" then SHout <= '1' after delay1 + 207*delay_incr;
elsif nramp = '0' and StoredData = "000011010000" then SHout <= '1' after delay1 + 208*delay_incr;
elsif nramp = '0' and StoredData = "000011010001" then SHout <= '1' after delay1 + 209*delay_incr;
elsif nramp = '0' and StoredData = "000011010010" then SHout <= '1' after delay1 + 210*delay_incr;
elsif nramp = '0' and StoredData = "000011010011" then SHout <= '1' after delay1 + 211*delay_incr;
elsif nramp = '0' and StoredData = "000011010100" then SHout <= '1' after delay1 + 212*delay_incr;
elsif nramp = '0' and StoredData = "000011010101" then SHout <= '1' after delay1 + 213*delay_incr;
elsif nramp = '0' and StoredData = "000011010110" then SHout <= '1' after delay1 + 214*delay_incr;
elsif nramp = '0' and StoredData = "000011010111" then SHout <= '1' after delay1 + 215*delay_incr;
elsif nramp = '0' and StoredData = "000011011000" then SHout <= '1' after delay1 + 216*delay_incr;
elsif nramp = '0' and StoredData = "000011011001" then SHout <= '1' after delay1 + 217*delay_incr;
elsif nramp = '0' and StoredData = "000011011010" then SHout <= '1' after delay1 + 218*delay_incr;
elsif nramp = '0' and StoredData = "000011011011" then SHout <= '1' after delay1 + 219*delay_incr;
elsif nramp = '0' and StoredData = "000011011100" then SHout <= '1' after delay1 + 220*delay_incr;
elsif nramp = '0' and StoredData = "000011011101" then SHout <= '1' after delay1 + 221*delay_incr;
elsif nramp = '0' and StoredData = "000011011110" then SHout <= '1' after delay1 + 222*delay_incr;
elsif nramp = '0' and StoredData = "000011011111" then SHout <= '1' after delay1 + 223*delay_incr;
elsif nramp = '0' and StoredData = "000011100000" then SHout <= '1' after delay1 + 224*delay_incr;
elsif nramp = '0' and StoredData = "000011100001" then SHout <= '1' after delay1 + 225*delay_incr;
elsif nramp = '0' and StoredData = "000011100010" then SHout <= '1' after delay1 + 226*delay_incr;
elsif nramp = '0' and StoredData = "000011100011" then SHout <= '1' after delay1 + 227*delay_incr;
elsif nramp = '0' and StoredData = "000011100100" then SHout <= '1' after delay1 + 228*delay_incr;
elsif nramp = '0' and StoredData = "000011100101" then SHout <= '1' after delay1 + 229*delay_incr;
elsif nramp = '0' and StoredData = "000011100110" then SHout <= '1' after delay1 + 230*delay_incr;
elsif nramp = '0' and StoredData = "000011100111" then SHout <= '1' after delay1 + 231*delay_incr;
elsif nramp = '0' and StoredData = "000011101000" then SHout <= '1' after delay1 + 232*delay_incr;
elsif nramp = '0' and StoredData = "000011101001" then SHout <= '1' after delay1 + 233*delay_incr;
elsif nramp = '0' and StoredData = "000011101010" then SHout <= '1' after delay1 + 234*delay_incr;
elsif nramp = '0' and StoredData = "000011101011" then SHout <= '1' after delay1 + 235*delay_incr;
elsif nramp = '0' and StoredData = "000011101100" then SHout <= '1' after delay1 + 236*delay_incr;
elsif nramp = '0' and StoredData = "000011101101" then SHout <= '1' after delay1 + 237*delay_incr;
elsif nramp = '0' and StoredData = "000011101110" then SHout <= '1' after delay1 + 238*delay_incr;
elsif nramp = '0' and StoredData = "000011101111" then SHout <= '1' after delay1 + 239*delay_incr;
elsif nramp = '0' and StoredData = "000011110000" then SHout <= '1' after delay1 + 240*delay_incr;
elsif nramp = '0' and StoredData = "000011110001" then SHout <= '1' after delay1 + 241*delay_incr;
elsif nramp = '0' and StoredData = "000011110010" then SHout <= '1' after delay1 + 242*delay_incr;
elsif nramp = '0' and StoredData = "000011110011" then SHout <= '1' after delay1 + 243*delay_incr;
elsif nramp = '0' and StoredData = "000011110100" then SHout <= '1' after delay1 + 244*delay_incr;
elsif nramp = '0' and StoredData = "000011110101" then SHout <= '1' after delay1 + 245*delay_incr;
elsif nramp = '0' and StoredData = "000011110110" then SHout <= '1' after delay1 + 246*delay_incr;
elsif nramp = '0' and StoredData = "000011110111" then SHout <= '1' after delay1 + 247*delay_incr;
elsif nramp = '0' and StoredData = "000011111000" then SHout <= '1' after delay1 + 248*delay_incr;
elsif nramp = '0' and StoredData = "000011111001" then SHout <= '1' after delay1 + 249*delay_incr;
elsif nramp = '0' and StoredData = "000011111010" then SHout <= '1' after delay1 + 250*delay_incr;
elsif nramp = '0' and StoredData = "000011111011" then SHout <= '1' after delay1 + 251*delay_incr;
elsif nramp = '0' and StoredData = "000011111100" then SHout <= '1' after delay1 + 252*delay_incr;
elsif nramp = '0' and StoredData = "000011111101" then SHout <= '1' after delay1 + 253*delay_incr;
elsif nramp = '0' and StoredData = "000011111110" then SHout <= '1' after delay1 + 254*delay_incr;
elsif nramp = '0' and StoredData = "000011111111" then SHout <= '1' after delay1 + 255*delay_incr;
elsif nramp = '0' and StoredData = "000100000000" then SHout <= '1' after delay1 + 256*delay_incr;
elsif nramp = '0' and StoredData = "000100000001" then SHout <= '1' after delay1 + 257*delay_incr;
elsif nramp = '0' and StoredData = "000100000010" then SHout <= '1' after delay1 + 258*delay_incr;
elsif nramp = '0' and StoredData = "000100000011" then SHout <= '1' after delay1 + 259*delay_incr;
elsif nramp = '0' and StoredData = "000100000100" then SHout <= '1' after delay1 + 260*delay_incr;
elsif nramp = '0' and StoredData = "000100000101" then SHout <= '1' after delay1 + 261*delay_incr;
elsif nramp = '0' and StoredData = "000100000110" then SHout <= '1' after delay1 + 262*delay_incr;
elsif nramp = '0' and StoredData = "000100000111" then SHout <= '1' after delay1 + 263*delay_incr;
elsif nramp = '0' and StoredData = "000100001000" then SHout <= '1' after delay1 + 264*delay_incr;
elsif nramp = '0' and StoredData = "000100001001" then SHout <= '1' after delay1 + 265*delay_incr;
elsif nramp = '0' and StoredData = "000100001010" then SHout <= '1' after delay1 + 266*delay_incr;
elsif nramp = '0' and StoredData = "000100001011" then SHout <= '1' after delay1 + 267*delay_incr;
elsif nramp = '0' and StoredData = "000100001100" then SHout <= '1' after delay1 + 268*delay_incr;
elsif nramp = '0' and StoredData = "000100001101" then SHout <= '1' after delay1 + 269*delay_incr;
elsif nramp = '0' and StoredData = "000100001110" then SHout <= '1' after delay1 + 270*delay_incr;
elsif nramp = '0' and StoredData = "000100001111" then SHout <= '1' after delay1 + 271*delay_incr;
elsif nramp = '0' and StoredData = "000100010000" then SHout <= '1' after delay1 + 272*delay_incr;
elsif nramp = '0' and StoredData = "000100010001" then SHout <= '1' after delay1 + 273*delay_incr;
elsif nramp = '0' and StoredData = "000100010010" then SHout <= '1' after delay1 + 274*delay_incr;
elsif nramp = '0' and StoredData = "000100010011" then SHout <= '1' after delay1 + 275*delay_incr;
elsif nramp = '0' and StoredData = "000100010100" then SHout <= '1' after delay1 + 276*delay_incr;
elsif nramp = '0' and StoredData = "000100010101" then SHout <= '1' after delay1 + 277*delay_incr;
elsif nramp = '0' and StoredData = "000100010110" then SHout <= '1' after delay1 + 278*delay_incr;
elsif nramp = '0' and StoredData = "000100010111" then SHout <= '1' after delay1 + 279*delay_incr;
elsif nramp = '0' and StoredData = "000100011000" then SHout <= '1' after delay1 + 280*delay_incr;
elsif nramp = '0' and StoredData = "000100011001" then SHout <= '1' after delay1 + 281*delay_incr;
elsif nramp = '0' and StoredData = "000100011010" then SHout <= '1' after delay1 + 282*delay_incr;
elsif nramp = '0' and StoredData = "000100011011" then SHout <= '1' after delay1 + 283*delay_incr;
elsif nramp = '0' and StoredData = "000100011100" then SHout <= '1' after delay1 + 284*delay_incr;
elsif nramp = '0' and StoredData = "000100011101" then SHout <= '1' after delay1 + 285*delay_incr;
elsif nramp = '0' and StoredData = "000100011110" then SHout <= '1' after delay1 + 286*delay_incr;
elsif nramp = '0' and StoredData = "000100011111" then SHout <= '1' after delay1 + 287*delay_incr;
elsif nramp = '0' and StoredData = "000100100000" then SHout <= '1' after delay1 + 288*delay_incr;
elsif nramp = '0' and StoredData = "000100100001" then SHout <= '1' after delay1 + 289*delay_incr;
elsif nramp = '0' and StoredData = "000100100010" then SHout <= '1' after delay1 + 290*delay_incr;
elsif nramp = '0' and StoredData = "000100100011" then SHout <= '1' after delay1 + 291*delay_incr;
elsif nramp = '0' and StoredData = "000100100100" then SHout <= '1' after delay1 + 292*delay_incr;
elsif nramp = '0' and StoredData = "000100100101" then SHout <= '1' after delay1 + 293*delay_incr;
elsif nramp = '0' and StoredData = "000100100110" then SHout <= '1' after delay1 + 294*delay_incr;
elsif nramp = '0' and StoredData = "000100100111" then SHout <= '1' after delay1 + 295*delay_incr;
elsif nramp = '0' and StoredData = "000100101000" then SHout <= '1' after delay1 + 296*delay_incr;
elsif nramp = '0' and StoredData = "000100101001" then SHout <= '1' after delay1 + 297*delay_incr;
elsif nramp = '0' and StoredData = "000100101010" then SHout <= '1' after delay1 + 298*delay_incr;
elsif nramp = '0' and StoredData = "000100101011" then SHout <= '1' after delay1 + 299*delay_incr;
elsif nramp = '0' and StoredData = "000100101100" then SHout <= '1' after delay1 + 300*delay_incr;
elsif nramp = '0' and StoredData = "000100101101" then SHout <= '1' after delay1 + 301*delay_incr;
elsif nramp = '0' and StoredData = "000100101110" then SHout <= '1' after delay1 + 302*delay_incr;
elsif nramp = '0' and StoredData = "000100101111" then SHout <= '1' after delay1 + 303*delay_incr;
elsif nramp = '0' and StoredData = "000100110000" then SHout <= '1' after delay1 + 304*delay_incr;
elsif nramp = '0' and StoredData = "000100110001" then SHout <= '1' after delay1 + 305*delay_incr;
elsif nramp = '0' and StoredData = "000100110010" then SHout <= '1' after delay1 + 306*delay_incr;
elsif nramp = '0' and StoredData = "000100110011" then SHout <= '1' after delay1 + 307*delay_incr;
elsif nramp = '0' and StoredData = "000100110100" then SHout <= '1' after delay1 + 308*delay_incr;
elsif nramp = '0' and StoredData = "000100110101" then SHout <= '1' after delay1 + 309*delay_incr;
elsif nramp = '0' and StoredData = "000100110110" then SHout <= '1' after delay1 + 310*delay_incr;
elsif nramp = '0' and StoredData = "000100110111" then SHout <= '1' after delay1 + 311*delay_incr;
elsif nramp = '0' and StoredData = "000100111000" then SHout <= '1' after delay1 + 312*delay_incr;
elsif nramp = '0' and StoredData = "000100111001" then SHout <= '1' after delay1 + 313*delay_incr;
elsif nramp = '0' and StoredData = "000100111010" then SHout <= '1' after delay1 + 314*delay_incr;
elsif nramp = '0' and StoredData = "000100111011" then SHout <= '1' after delay1 + 315*delay_incr;
elsif nramp = '0' and StoredData = "000100111100" then SHout <= '1' after delay1 + 316*delay_incr;
elsif nramp = '0' and StoredData = "000100111101" then SHout <= '1' after delay1 + 317*delay_incr;
elsif nramp = '0' and StoredData = "000100111110" then SHout <= '1' after delay1 + 318*delay_incr;
elsif nramp = '0' and StoredData = "000100111111" then SHout <= '1' after delay1 + 319*delay_incr;
elsif nramp = '0' and StoredData = "000101000000" then SHout <= '1' after delay1 + 320*delay_incr;
elsif nramp = '0' and StoredData = "000101000001" then SHout <= '1' after delay1 + 321*delay_incr;
elsif nramp = '0' and StoredData = "000101000010" then SHout <= '1' after delay1 + 322*delay_incr;
elsif nramp = '0' and StoredData = "000101000011" then SHout <= '1' after delay1 + 323*delay_incr;
elsif nramp = '0' and StoredData = "000101000100" then SHout <= '1' after delay1 + 324*delay_incr;
elsif nramp = '0' and StoredData = "000101000101" then SHout <= '1' after delay1 + 325*delay_incr;
elsif nramp = '0' and StoredData = "000101000110" then SHout <= '1' after delay1 + 326*delay_incr;
elsif nramp = '0' and StoredData = "000101000111" then SHout <= '1' after delay1 + 327*delay_incr;
elsif nramp = '0' and StoredData = "000101001000" then SHout <= '1' after delay1 + 328*delay_incr;
elsif nramp = '0' and StoredData = "000101001001" then SHout <= '1' after delay1 + 329*delay_incr;
elsif nramp = '0' and StoredData = "000101001010" then SHout <= '1' after delay1 + 330*delay_incr;
elsif nramp = '0' and StoredData = "000101001011" then SHout <= '1' after delay1 + 331*delay_incr;
elsif nramp = '0' and StoredData = "000101001100" then SHout <= '1' after delay1 + 332*delay_incr;
elsif nramp = '0' and StoredData = "000101001101" then SHout <= '1' after delay1 + 333*delay_incr;
elsif nramp = '0' and StoredData = "000101001110" then SHout <= '1' after delay1 + 334*delay_incr;
elsif nramp = '0' and StoredData = "000101001111" then SHout <= '1' after delay1 + 335*delay_incr;
elsif nramp = '0' and StoredData = "000101010000" then SHout <= '1' after delay1 + 336*delay_incr;
elsif nramp = '0' and StoredData = "000101010001" then SHout <= '1' after delay1 + 337*delay_incr;
elsif nramp = '0' and StoredData = "000101010010" then SHout <= '1' after delay1 + 338*delay_incr;
elsif nramp = '0' and StoredData = "000101010011" then SHout <= '1' after delay1 + 339*delay_incr;
elsif nramp = '0' and StoredData = "000101010100" then SHout <= '1' after delay1 + 340*delay_incr;
elsif nramp = '0' and StoredData = "000101010101" then SHout <= '1' after delay1 + 341*delay_incr;
elsif nramp = '0' and StoredData = "000101010110" then SHout <= '1' after delay1 + 342*delay_incr;
elsif nramp = '0' and StoredData = "000101010111" then SHout <= '1' after delay1 + 343*delay_incr;
elsif nramp = '0' and StoredData = "000101011000" then SHout <= '1' after delay1 + 344*delay_incr;
elsif nramp = '0' and StoredData = "000101011001" then SHout <= '1' after delay1 + 345*delay_incr;
elsif nramp = '0' and StoredData = "000101011010" then SHout <= '1' after delay1 + 346*delay_incr;
elsif nramp = '0' and StoredData = "000101011011" then SHout <= '1' after delay1 + 347*delay_incr;
elsif nramp = '0' and StoredData = "000101011100" then SHout <= '1' after delay1 + 348*delay_incr;
elsif nramp = '0' and StoredData = "000101011101" then SHout <= '1' after delay1 + 349*delay_incr;
elsif nramp = '0' and StoredData = "000101011110" then SHout <= '1' after delay1 + 350*delay_incr;
elsif nramp = '0' and StoredData = "000101011111" then SHout <= '1' after delay1 + 351*delay_incr;
elsif nramp = '0' and StoredData = "000101100000" then SHout <= '1' after delay1 + 352*delay_incr;
elsif nramp = '0' and StoredData = "000101100001" then SHout <= '1' after delay1 + 353*delay_incr;
elsif nramp = '0' and StoredData = "000101100010" then SHout <= '1' after delay1 + 354*delay_incr;
elsif nramp = '0' and StoredData = "000101100011" then SHout <= '1' after delay1 + 355*delay_incr;
elsif nramp = '0' and StoredData = "000101100100" then SHout <= '1' after delay1 + 356*delay_incr;
elsif nramp = '0' and StoredData = "000101100101" then SHout <= '1' after delay1 + 357*delay_incr;
elsif nramp = '0' and StoredData = "000101100110" then SHout <= '1' after delay1 + 358*delay_incr;
elsif nramp = '0' and StoredData = "000101100111" then SHout <= '1' after delay1 + 359*delay_incr;
elsif nramp = '0' and StoredData = "000101101000" then SHout <= '1' after delay1 + 360*delay_incr;
elsif nramp = '0' and StoredData = "000101101001" then SHout <= '1' after delay1 + 361*delay_incr;
elsif nramp = '0' and StoredData = "000101101010" then SHout <= '1' after delay1 + 362*delay_incr;
elsif nramp = '0' and StoredData = "000101101011" then SHout <= '1' after delay1 + 363*delay_incr;
elsif nramp = '0' and StoredData = "000101101100" then SHout <= '1' after delay1 + 364*delay_incr;
elsif nramp = '0' and StoredData = "000101101101" then SHout <= '1' after delay1 + 365*delay_incr;
elsif nramp = '0' and StoredData = "000101101110" then SHout <= '1' after delay1 + 366*delay_incr;
elsif nramp = '0' and StoredData = "000101101111" then SHout <= '1' after delay1 + 367*delay_incr;
elsif nramp = '0' and StoredData = "000101110000" then SHout <= '1' after delay1 + 368*delay_incr;
elsif nramp = '0' and StoredData = "000101110001" then SHout <= '1' after delay1 + 369*delay_incr;
elsif nramp = '0' and StoredData = "000101110010" then SHout <= '1' after delay1 + 370*delay_incr;
elsif nramp = '0' and StoredData = "000101110011" then SHout <= '1' after delay1 + 371*delay_incr;
elsif nramp = '0' and StoredData = "000101110100" then SHout <= '1' after delay1 + 372*delay_incr;
elsif nramp = '0' and StoredData = "000101110101" then SHout <= '1' after delay1 + 373*delay_incr;
elsif nramp = '0' and StoredData = "000101110110" then SHout <= '1' after delay1 + 374*delay_incr;
elsif nramp = '0' and StoredData = "000101110111" then SHout <= '1' after delay1 + 375*delay_incr;
elsif nramp = '0' and StoredData = "000101111000" then SHout <= '1' after delay1 + 376*delay_incr;
elsif nramp = '0' and StoredData = "000101111001" then SHout <= '1' after delay1 + 377*delay_incr;
elsif nramp = '0' and StoredData = "000101111010" then SHout <= '1' after delay1 + 378*delay_incr;
elsif nramp = '0' and StoredData = "000101111011" then SHout <= '1' after delay1 + 379*delay_incr;
elsif nramp = '0' and StoredData = "000101111100" then SHout <= '1' after delay1 + 380*delay_incr;
elsif nramp = '0' and StoredData = "000101111101" then SHout <= '1' after delay1 + 381*delay_incr;
elsif nramp = '0' and StoredData = "000101111110" then SHout <= '1' after delay1 + 382*delay_incr;
elsif nramp = '0' and StoredData = "000101111111" then SHout <= '1' after delay1 + 383*delay_incr;
elsif nramp = '0' and StoredData = "000110000000" then SHout <= '1' after delay1 + 384*delay_incr;
elsif nramp = '0' and StoredData = "000110000001" then SHout <= '1' after delay1 + 385*delay_incr;
elsif nramp = '0' and StoredData = "000110000010" then SHout <= '1' after delay1 + 386*delay_incr;
elsif nramp = '0' and StoredData = "000110000011" then SHout <= '1' after delay1 + 387*delay_incr;
elsif nramp = '0' and StoredData = "000110000100" then SHout <= '1' after delay1 + 388*delay_incr;
elsif nramp = '0' and StoredData = "000110000101" then SHout <= '1' after delay1 + 389*delay_incr;
elsif nramp = '0' and StoredData = "000110000110" then SHout <= '1' after delay1 + 390*delay_incr;
elsif nramp = '0' and StoredData = "000110000111" then SHout <= '1' after delay1 + 391*delay_incr;
elsif nramp = '0' and StoredData = "000110001000" then SHout <= '1' after delay1 + 392*delay_incr;
elsif nramp = '0' and StoredData = "000110001001" then SHout <= '1' after delay1 + 393*delay_incr;
elsif nramp = '0' and StoredData = "000110001010" then SHout <= '1' after delay1 + 394*delay_incr;
elsif nramp = '0' and StoredData = "000110001011" then SHout <= '1' after delay1 + 395*delay_incr;
elsif nramp = '0' and StoredData = "000110001100" then SHout <= '1' after delay1 + 396*delay_incr;
elsif nramp = '0' and StoredData = "000110001101" then SHout <= '1' after delay1 + 397*delay_incr;
elsif nramp = '0' and StoredData = "000110001110" then SHout <= '1' after delay1 + 398*delay_incr;
elsif nramp = '0' and StoredData = "000110001111" then SHout <= '1' after delay1 + 399*delay_incr;
elsif nramp = '0' and StoredData = "000110010000" then SHout <= '1' after delay1 + 400*delay_incr;
elsif nramp = '0' and StoredData = "000110010001" then SHout <= '1' after delay1 + 401*delay_incr;
elsif nramp = '0' and StoredData = "000110010010" then SHout <= '1' after delay1 + 402*delay_incr;
elsif nramp = '0' and StoredData = "000110010011" then SHout <= '1' after delay1 + 403*delay_incr;
elsif nramp = '0' and StoredData = "000110010100" then SHout <= '1' after delay1 + 404*delay_incr;
elsif nramp = '0' and StoredData = "000110010101" then SHout <= '1' after delay1 + 405*delay_incr;
elsif nramp = '0' and StoredData = "000110010110" then SHout <= '1' after delay1 + 406*delay_incr;
elsif nramp = '0' and StoredData = "000110010111" then SHout <= '1' after delay1 + 407*delay_incr;
elsif nramp = '0' and StoredData = "000110011000" then SHout <= '1' after delay1 + 408*delay_incr;
elsif nramp = '0' and StoredData = "000110011001" then SHout <= '1' after delay1 + 409*delay_incr;
elsif nramp = '0' and StoredData = "000110011010" then SHout <= '1' after delay1 + 410*delay_incr;
elsif nramp = '0' and StoredData = "000110011011" then SHout <= '1' after delay1 + 411*delay_incr;
elsif nramp = '0' and StoredData = "000110011100" then SHout <= '1' after delay1 + 412*delay_incr;
elsif nramp = '0' and StoredData = "000110011101" then SHout <= '1' after delay1 + 413*delay_incr;
elsif nramp = '0' and StoredData = "000110011110" then SHout <= '1' after delay1 + 414*delay_incr;
elsif nramp = '0' and StoredData = "000110011111" then SHout <= '1' after delay1 + 415*delay_incr;
elsif nramp = '0' and StoredData = "000110100000" then SHout <= '1' after delay1 + 416*delay_incr;
elsif nramp = '0' and StoredData = "000110100001" then SHout <= '1' after delay1 + 417*delay_incr;
elsif nramp = '0' and StoredData = "000110100010" then SHout <= '1' after delay1 + 418*delay_incr;
elsif nramp = '0' and StoredData = "000110100011" then SHout <= '1' after delay1 + 419*delay_incr;
elsif nramp = '0' and StoredData = "000110100100" then SHout <= '1' after delay1 + 420*delay_incr;
elsif nramp = '0' and StoredData = "000110100101" then SHout <= '1' after delay1 + 421*delay_incr;
elsif nramp = '0' and StoredData = "000110100110" then SHout <= '1' after delay1 + 422*delay_incr;
elsif nramp = '0' and StoredData = "000110100111" then SHout <= '1' after delay1 + 423*delay_incr;
elsif nramp = '0' and StoredData = "000110101000" then SHout <= '1' after delay1 + 424*delay_incr;
elsif nramp = '0' and StoredData = "000110101001" then SHout <= '1' after delay1 + 425*delay_incr;
elsif nramp = '0' and StoredData = "000110101010" then SHout <= '1' after delay1 + 426*delay_incr;
elsif nramp = '0' and StoredData = "000110101011" then SHout <= '1' after delay1 + 427*delay_incr;
elsif nramp = '0' and StoredData = "000110101100" then SHout <= '1' after delay1 + 428*delay_incr;
elsif nramp = '0' and StoredData = "000110101101" then SHout <= '1' after delay1 + 429*delay_incr;
elsif nramp = '0' and StoredData = "000110101110" then SHout <= '1' after delay1 + 430*delay_incr;
elsif nramp = '0' and StoredData = "000110101111" then SHout <= '1' after delay1 + 431*delay_incr;
elsif nramp = '0' and StoredData = "000110110000" then SHout <= '1' after delay1 + 432*delay_incr;
elsif nramp = '0' and StoredData = "000110110001" then SHout <= '1' after delay1 + 433*delay_incr;
elsif nramp = '0' and StoredData = "000110110010" then SHout <= '1' after delay1 + 434*delay_incr;
elsif nramp = '0' and StoredData = "000110110011" then SHout <= '1' after delay1 + 435*delay_incr;
elsif nramp = '0' and StoredData = "000110110100" then SHout <= '1' after delay1 + 436*delay_incr;
elsif nramp = '0' and StoredData = "000110110101" then SHout <= '1' after delay1 + 437*delay_incr;
elsif nramp = '0' and StoredData = "000110110110" then SHout <= '1' after delay1 + 438*delay_incr;
elsif nramp = '0' and StoredData = "000110110111" then SHout <= '1' after delay1 + 439*delay_incr;
elsif nramp = '0' and StoredData = "000110111000" then SHout <= '1' after delay1 + 440*delay_incr;
elsif nramp = '0' and StoredData = "000110111001" then SHout <= '1' after delay1 + 441*delay_incr;
elsif nramp = '0' and StoredData = "000110111010" then SHout <= '1' after delay1 + 442*delay_incr;
elsif nramp = '0' and StoredData = "000110111011" then SHout <= '1' after delay1 + 443*delay_incr;
elsif nramp = '0' and StoredData = "000110111100" then SHout <= '1' after delay1 + 444*delay_incr;
elsif nramp = '0' and StoredData = "000110111101" then SHout <= '1' after delay1 + 445*delay_incr;
elsif nramp = '0' and StoredData = "000110111110" then SHout <= '1' after delay1 + 446*delay_incr;
elsif nramp = '0' and StoredData = "000110111111" then SHout <= '1' after delay1 + 447*delay_incr;
elsif nramp = '0' and StoredData = "000111000000" then SHout <= '1' after delay1 + 448*delay_incr;
elsif nramp = '0' and StoredData = "000111000001" then SHout <= '1' after delay1 + 449*delay_incr;
elsif nramp = '0' and StoredData = "000111000010" then SHout <= '1' after delay1 + 450*delay_incr;
elsif nramp = '0' and StoredData = "000111000011" then SHout <= '1' after delay1 + 451*delay_incr;
elsif nramp = '0' and StoredData = "000111000100" then SHout <= '1' after delay1 + 452*delay_incr;
elsif nramp = '0' and StoredData = "000111000101" then SHout <= '1' after delay1 + 453*delay_incr;
elsif nramp = '0' and StoredData = "000111000110" then SHout <= '1' after delay1 + 454*delay_incr;
elsif nramp = '0' and StoredData = "000111000111" then SHout <= '1' after delay1 + 455*delay_incr;
elsif nramp = '0' and StoredData = "000111001000" then SHout <= '1' after delay1 + 456*delay_incr;
elsif nramp = '0' and StoredData = "000111001001" then SHout <= '1' after delay1 + 457*delay_incr;
elsif nramp = '0' and StoredData = "000111001010" then SHout <= '1' after delay1 + 458*delay_incr;
elsif nramp = '0' and StoredData = "000111001011" then SHout <= '1' after delay1 + 459*delay_incr;
elsif nramp = '0' and StoredData = "000111001100" then SHout <= '1' after delay1 + 460*delay_incr;
elsif nramp = '0' and StoredData = "000111001101" then SHout <= '1' after delay1 + 461*delay_incr;
elsif nramp = '0' and StoredData = "000111001110" then SHout <= '1' after delay1 + 462*delay_incr;
elsif nramp = '0' and StoredData = "000111001111" then SHout <= '1' after delay1 + 463*delay_incr;
elsif nramp = '0' and StoredData = "000111010000" then SHout <= '1' after delay1 + 464*delay_incr;
elsif nramp = '0' and StoredData = "000111010001" then SHout <= '1' after delay1 + 465*delay_incr;
elsif nramp = '0' and StoredData = "000111010010" then SHout <= '1' after delay1 + 466*delay_incr;
elsif nramp = '0' and StoredData = "000111010011" then SHout <= '1' after delay1 + 467*delay_incr;
elsif nramp = '0' and StoredData = "000111010100" then SHout <= '1' after delay1 + 468*delay_incr;
elsif nramp = '0' and StoredData = "000111010101" then SHout <= '1' after delay1 + 469*delay_incr;
elsif nramp = '0' and StoredData = "000111010110" then SHout <= '1' after delay1 + 470*delay_incr;
elsif nramp = '0' and StoredData = "000111010111" then SHout <= '1' after delay1 + 471*delay_incr;
elsif nramp = '0' and StoredData = "000111011000" then SHout <= '1' after delay1 + 472*delay_incr;
elsif nramp = '0' and StoredData = "000111011001" then SHout <= '1' after delay1 + 473*delay_incr;
elsif nramp = '0' and StoredData = "000111011010" then SHout <= '1' after delay1 + 474*delay_incr;
elsif nramp = '0' and StoredData = "000111011011" then SHout <= '1' after delay1 + 475*delay_incr;
elsif nramp = '0' and StoredData = "000111011100" then SHout <= '1' after delay1 + 476*delay_incr;
elsif nramp = '0' and StoredData = "000111011101" then SHout <= '1' after delay1 + 477*delay_incr;
elsif nramp = '0' and StoredData = "000111011110" then SHout <= '1' after delay1 + 478*delay_incr;
elsif nramp = '0' and StoredData = "000111011111" then SHout <= '1' after delay1 + 479*delay_incr;
elsif nramp = '0' and StoredData = "000111100000" then SHout <= '1' after delay1 + 480*delay_incr;
elsif nramp = '0' and StoredData = "000111100001" then SHout <= '1' after delay1 + 481*delay_incr;
elsif nramp = '0' and StoredData = "000111100010" then SHout <= '1' after delay1 + 482*delay_incr;
elsif nramp = '0' and StoredData = "000111100011" then SHout <= '1' after delay1 + 483*delay_incr;
elsif nramp = '0' and StoredData = "000111100100" then SHout <= '1' after delay1 + 484*delay_incr;
elsif nramp = '0' and StoredData = "000111100101" then SHout <= '1' after delay1 + 485*delay_incr;
elsif nramp = '0' and StoredData = "000111100110" then SHout <= '1' after delay1 + 486*delay_incr;
elsif nramp = '0' and StoredData = "000111100111" then SHout <= '1' after delay1 + 487*delay_incr;
elsif nramp = '0' and StoredData = "000111101000" then SHout <= '1' after delay1 + 488*delay_incr;
elsif nramp = '0' and StoredData = "000111101001" then SHout <= '1' after delay1 + 489*delay_incr;
elsif nramp = '0' and StoredData = "000111101010" then SHout <= '1' after delay1 + 490*delay_incr;
elsif nramp = '0' and StoredData = "000111101011" then SHout <= '1' after delay1 + 491*delay_incr;
elsif nramp = '0' and StoredData = "000111101100" then SHout <= '1' after delay1 + 492*delay_incr;
elsif nramp = '0' and StoredData = "000111101101" then SHout <= '1' after delay1 + 493*delay_incr;
elsif nramp = '0' and StoredData = "000111101110" then SHout <= '1' after delay1 + 494*delay_incr;
elsif nramp = '0' and StoredData = "000111101111" then SHout <= '1' after delay1 + 495*delay_incr;
elsif nramp = '0' and StoredData = "000111110000" then SHout <= '1' after delay1 + 496*delay_incr;
elsif nramp = '0' and StoredData = "000111110001" then SHout <= '1' after delay1 + 497*delay_incr;
elsif nramp = '0' and StoredData = "000111110010" then SHout <= '1' after delay1 + 498*delay_incr;
elsif nramp = '0' and StoredData = "000111110011" then SHout <= '1' after delay1 + 499*delay_incr;
elsif nramp = '0' and StoredData = "000111110100" then SHout <= '1' after delay1 + 500*delay_incr;
elsif nramp = '0' and StoredData = "000111110101" then SHout <= '1' after delay1 + 501*delay_incr;
elsif nramp = '0' and StoredData = "000111110110" then SHout <= '1' after delay1 + 502*delay_incr;
elsif nramp = '0' and StoredData = "000111110111" then SHout <= '1' after delay1 + 503*delay_incr;
elsif nramp = '0' and StoredData = "000111111000" then SHout <= '1' after delay1 + 504*delay_incr;
elsif nramp = '0' and StoredData = "000111111001" then SHout <= '1' after delay1 + 505*delay_incr;
elsif nramp = '0' and StoredData = "000111111010" then SHout <= '1' after delay1 + 506*delay_incr;
elsif nramp = '0' and StoredData = "000111111011" then SHout <= '1' after delay1 + 507*delay_incr;
elsif nramp = '0' and StoredData = "000111111100" then SHout <= '1' after delay1 + 508*delay_incr;
elsif nramp = '0' and StoredData = "000111111101" then SHout <= '1' after delay1 + 509*delay_incr;
elsif nramp = '0' and StoredData = "000111111110" then SHout <= '1' after delay1 + 510*delay_incr;
elsif nramp = '0' and StoredData = "000111111111" then SHout <= '1' after delay1 + 511*delay_incr;
elsif nramp = '0' and StoredData = "001000000000" then SHout <= '1' after delay1 + 512*delay_incr;
elsif nramp = '0' and StoredData = "001000000001" then SHout <= '1' after delay1 + 513*delay_incr;
elsif nramp = '0' and StoredData = "001000000010" then SHout <= '1' after delay1 + 514*delay_incr;
elsif nramp = '0' and StoredData = "001000000011" then SHout <= '1' after delay1 + 515*delay_incr;
elsif nramp = '0' and StoredData = "001000000100" then SHout <= '1' after delay1 + 516*delay_incr;
elsif nramp = '0' and StoredData = "001000000101" then SHout <= '1' after delay1 + 517*delay_incr;
elsif nramp = '0' and StoredData = "001000000110" then SHout <= '1' after delay1 + 518*delay_incr;
elsif nramp = '0' and StoredData = "001000000111" then SHout <= '1' after delay1 + 519*delay_incr;
elsif nramp = '0' and StoredData = "001000001000" then SHout <= '1' after delay1 + 520*delay_incr;
elsif nramp = '0' and StoredData = "001000001001" then SHout <= '1' after delay1 + 521*delay_incr;
elsif nramp = '0' and StoredData = "001000001010" then SHout <= '1' after delay1 + 522*delay_incr;
elsif nramp = '0' and StoredData = "001000001011" then SHout <= '1' after delay1 + 523*delay_incr;
elsif nramp = '0' and StoredData = "001000001100" then SHout <= '1' after delay1 + 524*delay_incr;
elsif nramp = '0' and StoredData = "001000001101" then SHout <= '1' after delay1 + 525*delay_incr;
elsif nramp = '0' and StoredData = "001000001110" then SHout <= '1' after delay1 + 526*delay_incr;
elsif nramp = '0' and StoredData = "001000001111" then SHout <= '1' after delay1 + 527*delay_incr;
elsif nramp = '0' and StoredData = "001000010000" then SHout <= '1' after delay1 + 528*delay_incr;
elsif nramp = '0' and StoredData = "001000010001" then SHout <= '1' after delay1 + 529*delay_incr;
elsif nramp = '0' and StoredData = "001000010010" then SHout <= '1' after delay1 + 530*delay_incr;
elsif nramp = '0' and StoredData = "001000010011" then SHout <= '1' after delay1 + 531*delay_incr;
elsif nramp = '0' and StoredData = "001000010100" then SHout <= '1' after delay1 + 532*delay_incr;
elsif nramp = '0' and StoredData = "001000010101" then SHout <= '1' after delay1 + 533*delay_incr;
elsif nramp = '0' and StoredData = "001000010110" then SHout <= '1' after delay1 + 534*delay_incr;
elsif nramp = '0' and StoredData = "001000010111" then SHout <= '1' after delay1 + 535*delay_incr;
elsif nramp = '0' and StoredData = "001000011000" then SHout <= '1' after delay1 + 536*delay_incr;
elsif nramp = '0' and StoredData = "001000011001" then SHout <= '1' after delay1 + 537*delay_incr;
elsif nramp = '0' and StoredData = "001000011010" then SHout <= '1' after delay1 + 538*delay_incr;
elsif nramp = '0' and StoredData = "001000011011" then SHout <= '1' after delay1 + 539*delay_incr;
elsif nramp = '0' and StoredData = "001000011100" then SHout <= '1' after delay1 + 540*delay_incr;
elsif nramp = '0' and StoredData = "001000011101" then SHout <= '1' after delay1 + 541*delay_incr;
elsif nramp = '0' and StoredData = "001000011110" then SHout <= '1' after delay1 + 542*delay_incr;
elsif nramp = '0' and StoredData = "001000011111" then SHout <= '1' after delay1 + 543*delay_incr;
elsif nramp = '0' and StoredData = "001000100000" then SHout <= '1' after delay1 + 544*delay_incr;
elsif nramp = '0' and StoredData = "001000100001" then SHout <= '1' after delay1 + 545*delay_incr;
elsif nramp = '0' and StoredData = "001000100010" then SHout <= '1' after delay1 + 546*delay_incr;
elsif nramp = '0' and StoredData = "001000100011" then SHout <= '1' after delay1 + 547*delay_incr;
elsif nramp = '0' and StoredData = "001000100100" then SHout <= '1' after delay1 + 548*delay_incr;
elsif nramp = '0' and StoredData = "001000100101" then SHout <= '1' after delay1 + 549*delay_incr;
elsif nramp = '0' and StoredData = "001000100110" then SHout <= '1' after delay1 + 550*delay_incr;
elsif nramp = '0' and StoredData = "001000100111" then SHout <= '1' after delay1 + 551*delay_incr;
elsif nramp = '0' and StoredData = "001000101000" then SHout <= '1' after delay1 + 552*delay_incr;
elsif nramp = '0' and StoredData = "001000101001" then SHout <= '1' after delay1 + 553*delay_incr;
elsif nramp = '0' and StoredData = "001000101010" then SHout <= '1' after delay1 + 554*delay_incr;
elsif nramp = '0' and StoredData = "001000101011" then SHout <= '1' after delay1 + 555*delay_incr;
elsif nramp = '0' and StoredData = "001000101100" then SHout <= '1' after delay1 + 556*delay_incr;
elsif nramp = '0' and StoredData = "001000101101" then SHout <= '1' after delay1 + 557*delay_incr;
elsif nramp = '0' and StoredData = "001000101110" then SHout <= '1' after delay1 + 558*delay_incr;
elsif nramp = '0' and StoredData = "001000101111" then SHout <= '1' after delay1 + 559*delay_incr;
elsif nramp = '0' and StoredData = "001000110000" then SHout <= '1' after delay1 + 560*delay_incr;
elsif nramp = '0' and StoredData = "001000110001" then SHout <= '1' after delay1 + 561*delay_incr;
elsif nramp = '0' and StoredData = "001000110010" then SHout <= '1' after delay1 + 562*delay_incr;
elsif nramp = '0' and StoredData = "001000110011" then SHout <= '1' after delay1 + 563*delay_incr;
elsif nramp = '0' and StoredData = "001000110100" then SHout <= '1' after delay1 + 564*delay_incr;
elsif nramp = '0' and StoredData = "001000110101" then SHout <= '1' after delay1 + 565*delay_incr;
elsif nramp = '0' and StoredData = "001000110110" then SHout <= '1' after delay1 + 566*delay_incr;
elsif nramp = '0' and StoredData = "001000110111" then SHout <= '1' after delay1 + 567*delay_incr;
elsif nramp = '0' and StoredData = "001000111000" then SHout <= '1' after delay1 + 568*delay_incr;
elsif nramp = '0' and StoredData = "001000111001" then SHout <= '1' after delay1 + 569*delay_incr;
elsif nramp = '0' and StoredData = "001000111010" then SHout <= '1' after delay1 + 570*delay_incr;
elsif nramp = '0' and StoredData = "001000111011" then SHout <= '1' after delay1 + 571*delay_incr;
elsif nramp = '0' and StoredData = "001000111100" then SHout <= '1' after delay1 + 572*delay_incr;
elsif nramp = '0' and StoredData = "001000111101" then SHout <= '1' after delay1 + 573*delay_incr;
elsif nramp = '0' and StoredData = "001000111110" then SHout <= '1' after delay1 + 574*delay_incr;
elsif nramp = '0' and StoredData = "001000111111" then SHout <= '1' after delay1 + 575*delay_incr;
elsif nramp = '0' and StoredData = "001001000000" then SHout <= '1' after delay1 + 576*delay_incr;
elsif nramp = '0' and StoredData = "001001000001" then SHout <= '1' after delay1 + 577*delay_incr;
elsif nramp = '0' and StoredData = "001001000010" then SHout <= '1' after delay1 + 578*delay_incr;
elsif nramp = '0' and StoredData = "001001000011" then SHout <= '1' after delay1 + 579*delay_incr;
elsif nramp = '0' and StoredData = "001001000100" then SHout <= '1' after delay1 + 580*delay_incr;
elsif nramp = '0' and StoredData = "001001000101" then SHout <= '1' after delay1 + 581*delay_incr;
elsif nramp = '0' and StoredData = "001001000110" then SHout <= '1' after delay1 + 582*delay_incr;
elsif nramp = '0' and StoredData = "001001000111" then SHout <= '1' after delay1 + 583*delay_incr;
elsif nramp = '0' and StoredData = "001001001000" then SHout <= '1' after delay1 + 584*delay_incr;
elsif nramp = '0' and StoredData = "001001001001" then SHout <= '1' after delay1 + 585*delay_incr;
elsif nramp = '0' and StoredData = "001001001010" then SHout <= '1' after delay1 + 586*delay_incr;
elsif nramp = '0' and StoredData = "001001001011" then SHout <= '1' after delay1 + 587*delay_incr;
elsif nramp = '0' and StoredData = "001001001100" then SHout <= '1' after delay1 + 588*delay_incr;
elsif nramp = '0' and StoredData = "001001001101" then SHout <= '1' after delay1 + 589*delay_incr;
elsif nramp = '0' and StoredData = "001001001110" then SHout <= '1' after delay1 + 590*delay_incr;
elsif nramp = '0' and StoredData = "001001001111" then SHout <= '1' after delay1 + 591*delay_incr;
elsif nramp = '0' and StoredData = "001001010000" then SHout <= '1' after delay1 + 592*delay_incr;
elsif nramp = '0' and StoredData = "001001010001" then SHout <= '1' after delay1 + 593*delay_incr;
elsif nramp = '0' and StoredData = "001001010010" then SHout <= '1' after delay1 + 594*delay_incr;
elsif nramp = '0' and StoredData = "001001010011" then SHout <= '1' after delay1 + 595*delay_incr;
elsif nramp = '0' and StoredData = "001001010100" then SHout <= '1' after delay1 + 596*delay_incr;
elsif nramp = '0' and StoredData = "001001010101" then SHout <= '1' after delay1 + 597*delay_incr;
elsif nramp = '0' and StoredData = "001001010110" then SHout <= '1' after delay1 + 598*delay_incr;
elsif nramp = '0' and StoredData = "001001010111" then SHout <= '1' after delay1 + 599*delay_incr;
elsif nramp = '0' and StoredData = "001001011000" then SHout <= '1' after delay1 + 600*delay_incr;
elsif nramp = '0' and StoredData = "001001011001" then SHout <= '1' after delay1 + 601*delay_incr;
elsif nramp = '0' and StoredData = "001001011010" then SHout <= '1' after delay1 + 602*delay_incr;
elsif nramp = '0' and StoredData = "001001011011" then SHout <= '1' after delay1 + 603*delay_incr;
elsif nramp = '0' and StoredData = "001001011100" then SHout <= '1' after delay1 + 604*delay_incr;
elsif nramp = '0' and StoredData = "001001011101" then SHout <= '1' after delay1 + 605*delay_incr;
elsif nramp = '0' and StoredData = "001001011110" then SHout <= '1' after delay1 + 606*delay_incr;
elsif nramp = '0' and StoredData = "001001011111" then SHout <= '1' after delay1 + 607*delay_incr;
elsif nramp = '0' and StoredData = "001001100000" then SHout <= '1' after delay1 + 608*delay_incr;
elsif nramp = '0' and StoredData = "001001100001" then SHout <= '1' after delay1 + 609*delay_incr;
elsif nramp = '0' and StoredData = "001001100010" then SHout <= '1' after delay1 + 610*delay_incr;
elsif nramp = '0' and StoredData = "001001100011" then SHout <= '1' after delay1 + 611*delay_incr;
elsif nramp = '0' and StoredData = "001001100100" then SHout <= '1' after delay1 + 612*delay_incr;
elsif nramp = '0' and StoredData = "001001100101" then SHout <= '1' after delay1 + 613*delay_incr;
elsif nramp = '0' and StoredData = "001001100110" then SHout <= '1' after delay1 + 614*delay_incr;
elsif nramp = '0' and StoredData = "001001100111" then SHout <= '1' after delay1 + 615*delay_incr;
elsif nramp = '0' and StoredData = "001001101000" then SHout <= '1' after delay1 + 616*delay_incr;
elsif nramp = '0' and StoredData = "001001101001" then SHout <= '1' after delay1 + 617*delay_incr;
elsif nramp = '0' and StoredData = "001001101010" then SHout <= '1' after delay1 + 618*delay_incr;
elsif nramp = '0' and StoredData = "001001101011" then SHout <= '1' after delay1 + 619*delay_incr;
elsif nramp = '0' and StoredData = "001001101100" then SHout <= '1' after delay1 + 620*delay_incr;
elsif nramp = '0' and StoredData = "001001101101" then SHout <= '1' after delay1 + 621*delay_incr;
elsif nramp = '0' and StoredData = "001001101110" then SHout <= '1' after delay1 + 622*delay_incr;
elsif nramp = '0' and StoredData = "001001101111" then SHout <= '1' after delay1 + 623*delay_incr;
elsif nramp = '0' and StoredData = "001001110000" then SHout <= '1' after delay1 + 624*delay_incr;
elsif nramp = '0' and StoredData = "001001110001" then SHout <= '1' after delay1 + 625*delay_incr;
elsif nramp = '0' and StoredData = "001001110010" then SHout <= '1' after delay1 + 626*delay_incr;
elsif nramp = '0' and StoredData = "001001110011" then SHout <= '1' after delay1 + 627*delay_incr;
elsif nramp = '0' and StoredData = "001001110100" then SHout <= '1' after delay1 + 628*delay_incr;
elsif nramp = '0' and StoredData = "001001110101" then SHout <= '1' after delay1 + 629*delay_incr;
elsif nramp = '0' and StoredData = "001001110110" then SHout <= '1' after delay1 + 630*delay_incr;
elsif nramp = '0' and StoredData = "001001110111" then SHout <= '1' after delay1 + 631*delay_incr;
elsif nramp = '0' and StoredData = "001001111000" then SHout <= '1' after delay1 + 632*delay_incr;
elsif nramp = '0' and StoredData = "001001111001" then SHout <= '1' after delay1 + 633*delay_incr;
elsif nramp = '0' and StoredData = "001001111010" then SHout <= '1' after delay1 + 634*delay_incr;
elsif nramp = '0' and StoredData = "001001111011" then SHout <= '1' after delay1 + 635*delay_incr;
elsif nramp = '0' and StoredData = "001001111100" then SHout <= '1' after delay1 + 636*delay_incr;
elsif nramp = '0' and StoredData = "001001111101" then SHout <= '1' after delay1 + 637*delay_incr;
elsif nramp = '0' and StoredData = "001001111110" then SHout <= '1' after delay1 + 638*delay_incr;
elsif nramp = '0' and StoredData = "001001111111" then SHout <= '1' after delay1 + 639*delay_incr;
elsif nramp = '0' and StoredData = "001010000000" then SHout <= '1' after delay1 + 640*delay_incr;
elsif nramp = '0' and StoredData = "001010000001" then SHout <= '1' after delay1 + 641*delay_incr;
elsif nramp = '0' and StoredData = "001010000010" then SHout <= '1' after delay1 + 642*delay_incr;
elsif nramp = '0' and StoredData = "001010000011" then SHout <= '1' after delay1 + 643*delay_incr;
elsif nramp = '0' and StoredData = "001010000100" then SHout <= '1' after delay1 + 644*delay_incr;
elsif nramp = '0' and StoredData = "001010000101" then SHout <= '1' after delay1 + 645*delay_incr;
elsif nramp = '0' and StoredData = "001010000110" then SHout <= '1' after delay1 + 646*delay_incr;
elsif nramp = '0' and StoredData = "001010000111" then SHout <= '1' after delay1 + 647*delay_incr;
elsif nramp = '0' and StoredData = "001010001000" then SHout <= '1' after delay1 + 648*delay_incr;
elsif nramp = '0' and StoredData = "001010001001" then SHout <= '1' after delay1 + 649*delay_incr;
elsif nramp = '0' and StoredData = "001010001010" then SHout <= '1' after delay1 + 650*delay_incr;
elsif nramp = '0' and StoredData = "001010001011" then SHout <= '1' after delay1 + 651*delay_incr;
elsif nramp = '0' and StoredData = "001010001100" then SHout <= '1' after delay1 + 652*delay_incr;
elsif nramp = '0' and StoredData = "001010001101" then SHout <= '1' after delay1 + 653*delay_incr;
elsif nramp = '0' and StoredData = "001010001110" then SHout <= '1' after delay1 + 654*delay_incr;
elsif nramp = '0' and StoredData = "001010001111" then SHout <= '1' after delay1 + 655*delay_incr;
elsif nramp = '0' and StoredData = "001010010000" then SHout <= '1' after delay1 + 656*delay_incr;
elsif nramp = '0' and StoredData = "001010010001" then SHout <= '1' after delay1 + 657*delay_incr;
elsif nramp = '0' and StoredData = "001010010010" then SHout <= '1' after delay1 + 658*delay_incr;
elsif nramp = '0' and StoredData = "001010010011" then SHout <= '1' after delay1 + 659*delay_incr;
elsif nramp = '0' and StoredData = "001010010100" then SHout <= '1' after delay1 + 660*delay_incr;
elsif nramp = '0' and StoredData = "001010010101" then SHout <= '1' after delay1 + 661*delay_incr;
elsif nramp = '0' and StoredData = "001010010110" then SHout <= '1' after delay1 + 662*delay_incr;
elsif nramp = '0' and StoredData = "001010010111" then SHout <= '1' after delay1 + 663*delay_incr;
elsif nramp = '0' and StoredData = "001010011000" then SHout <= '1' after delay1 + 664*delay_incr;
elsif nramp = '0' and StoredData = "001010011001" then SHout <= '1' after delay1 + 665*delay_incr;
elsif nramp = '0' and StoredData = "001010011010" then SHout <= '1' after delay1 + 666*delay_incr;
elsif nramp = '0' and StoredData = "001010011011" then SHout <= '1' after delay1 + 667*delay_incr;
elsif nramp = '0' and StoredData = "001010011100" then SHout <= '1' after delay1 + 668*delay_incr;
elsif nramp = '0' and StoredData = "001010011101" then SHout <= '1' after delay1 + 669*delay_incr;
elsif nramp = '0' and StoredData = "001010011110" then SHout <= '1' after delay1 + 670*delay_incr;
elsif nramp = '0' and StoredData = "001010011111" then SHout <= '1' after delay1 + 671*delay_incr;
elsif nramp = '0' and StoredData = "001010100000" then SHout <= '1' after delay1 + 672*delay_incr;
elsif nramp = '0' and StoredData = "001010100001" then SHout <= '1' after delay1 + 673*delay_incr;
elsif nramp = '0' and StoredData = "001010100010" then SHout <= '1' after delay1 + 674*delay_incr;
elsif nramp = '0' and StoredData = "001010100011" then SHout <= '1' after delay1 + 675*delay_incr;
elsif nramp = '0' and StoredData = "001010100100" then SHout <= '1' after delay1 + 676*delay_incr;
elsif nramp = '0' and StoredData = "001010100101" then SHout <= '1' after delay1 + 677*delay_incr;
elsif nramp = '0' and StoredData = "001010100110" then SHout <= '1' after delay1 + 678*delay_incr;
elsif nramp = '0' and StoredData = "001010100111" then SHout <= '1' after delay1 + 679*delay_incr;
elsif nramp = '0' and StoredData = "001010101000" then SHout <= '1' after delay1 + 680*delay_incr;
elsif nramp = '0' and StoredData = "001010101001" then SHout <= '1' after delay1 + 681*delay_incr;
elsif nramp = '0' and StoredData = "001010101010" then SHout <= '1' after delay1 + 682*delay_incr;
elsif nramp = '0' and StoredData = "001010101011" then SHout <= '1' after delay1 + 683*delay_incr;
elsif nramp = '0' and StoredData = "001010101100" then SHout <= '1' after delay1 + 684*delay_incr;
elsif nramp = '0' and StoredData = "001010101101" then SHout <= '1' after delay1 + 685*delay_incr;
elsif nramp = '0' and StoredData = "001010101110" then SHout <= '1' after delay1 + 686*delay_incr;
elsif nramp = '0' and StoredData = "001010101111" then SHout <= '1' after delay1 + 687*delay_incr;
elsif nramp = '0' and StoredData = "001010110000" then SHout <= '1' after delay1 + 688*delay_incr;
elsif nramp = '0' and StoredData = "001010110001" then SHout <= '1' after delay1 + 689*delay_incr;
elsif nramp = '0' and StoredData = "001010110010" then SHout <= '1' after delay1 + 690*delay_incr;
elsif nramp = '0' and StoredData = "001010110011" then SHout <= '1' after delay1 + 691*delay_incr;
elsif nramp = '0' and StoredData = "001010110100" then SHout <= '1' after delay1 + 692*delay_incr;
elsif nramp = '0' and StoredData = "001010110101" then SHout <= '1' after delay1 + 693*delay_incr;
elsif nramp = '0' and StoredData = "001010110110" then SHout <= '1' after delay1 + 694*delay_incr;
elsif nramp = '0' and StoredData = "001010110111" then SHout <= '1' after delay1 + 695*delay_incr;
elsif nramp = '0' and StoredData = "001010111000" then SHout <= '1' after delay1 + 696*delay_incr;
elsif nramp = '0' and StoredData = "001010111001" then SHout <= '1' after delay1 + 697*delay_incr;
elsif nramp = '0' and StoredData = "001010111010" then SHout <= '1' after delay1 + 698*delay_incr;
elsif nramp = '0' and StoredData = "001010111011" then SHout <= '1' after delay1 + 699*delay_incr;
elsif nramp = '0' and StoredData = "001010111100" then SHout <= '1' after delay1 + 700*delay_incr;
elsif nramp = '0' and StoredData = "001010111101" then SHout <= '1' after delay1 + 701*delay_incr;
elsif nramp = '0' and StoredData = "001010111110" then SHout <= '1' after delay1 + 702*delay_incr;
elsif nramp = '0' and StoredData = "001010111111" then SHout <= '1' after delay1 + 703*delay_incr;
elsif nramp = '0' and StoredData = "001011000000" then SHout <= '1' after delay1 + 704*delay_incr;
elsif nramp = '0' and StoredData = "001011000001" then SHout <= '1' after delay1 + 705*delay_incr;
elsif nramp = '0' and StoredData = "001011000010" then SHout <= '1' after delay1 + 706*delay_incr;
elsif nramp = '0' and StoredData = "001011000011" then SHout <= '1' after delay1 + 707*delay_incr;
elsif nramp = '0' and StoredData = "001011000100" then SHout <= '1' after delay1 + 708*delay_incr;
elsif nramp = '0' and StoredData = "001011000101" then SHout <= '1' after delay1 + 709*delay_incr;
elsif nramp = '0' and StoredData = "001011000110" then SHout <= '1' after delay1 + 710*delay_incr;
elsif nramp = '0' and StoredData = "001011000111" then SHout <= '1' after delay1 + 711*delay_incr;
elsif nramp = '0' and StoredData = "001011001000" then SHout <= '1' after delay1 + 712*delay_incr;
elsif nramp = '0' and StoredData = "001011001001" then SHout <= '1' after delay1 + 713*delay_incr;
elsif nramp = '0' and StoredData = "001011001010" then SHout <= '1' after delay1 + 714*delay_incr;
elsif nramp = '0' and StoredData = "001011001011" then SHout <= '1' after delay1 + 715*delay_incr;
elsif nramp = '0' and StoredData = "001011001100" then SHout <= '1' after delay1 + 716*delay_incr;
elsif nramp = '0' and StoredData = "001011001101" then SHout <= '1' after delay1 + 717*delay_incr;
elsif nramp = '0' and StoredData = "001011001110" then SHout <= '1' after delay1 + 718*delay_incr;
elsif nramp = '0' and StoredData = "001011001111" then SHout <= '1' after delay1 + 719*delay_incr;
elsif nramp = '0' and StoredData = "001011010000" then SHout <= '1' after delay1 + 720*delay_incr;
elsif nramp = '0' and StoredData = "001011010001" then SHout <= '1' after delay1 + 721*delay_incr;
elsif nramp = '0' and StoredData = "001011010010" then SHout <= '1' after delay1 + 722*delay_incr;
elsif nramp = '0' and StoredData = "001011010011" then SHout <= '1' after delay1 + 723*delay_incr;
elsif nramp = '0' and StoredData = "001011010100" then SHout <= '1' after delay1 + 724*delay_incr;
elsif nramp = '0' and StoredData = "001011010101" then SHout <= '1' after delay1 + 725*delay_incr;
elsif nramp = '0' and StoredData = "001011010110" then SHout <= '1' after delay1 + 726*delay_incr;
elsif nramp = '0' and StoredData = "001011010111" then SHout <= '1' after delay1 + 727*delay_incr;
elsif nramp = '0' and StoredData = "001011011000" then SHout <= '1' after delay1 + 728*delay_incr;
elsif nramp = '0' and StoredData = "001011011001" then SHout <= '1' after delay1 + 729*delay_incr;
elsif nramp = '0' and StoredData = "001011011010" then SHout <= '1' after delay1 + 730*delay_incr;
elsif nramp = '0' and StoredData = "001011011011" then SHout <= '1' after delay1 + 731*delay_incr;
elsif nramp = '0' and StoredData = "001011011100" then SHout <= '1' after delay1 + 732*delay_incr;
elsif nramp = '0' and StoredData = "001011011101" then SHout <= '1' after delay1 + 733*delay_incr;
elsif nramp = '0' and StoredData = "001011011110" then SHout <= '1' after delay1 + 734*delay_incr;
elsif nramp = '0' and StoredData = "001011011111" then SHout <= '1' after delay1 + 735*delay_incr;
elsif nramp = '0' and StoredData = "001011100000" then SHout <= '1' after delay1 + 736*delay_incr;
elsif nramp = '0' and StoredData = "001011100001" then SHout <= '1' after delay1 + 737*delay_incr;
elsif nramp = '0' and StoredData = "001011100010" then SHout <= '1' after delay1 + 738*delay_incr;
elsif nramp = '0' and StoredData = "001011100011" then SHout <= '1' after delay1 + 739*delay_incr;
elsif nramp = '0' and StoredData = "001011100100" then SHout <= '1' after delay1 + 740*delay_incr;
elsif nramp = '0' and StoredData = "001011100101" then SHout <= '1' after delay1 + 741*delay_incr;
elsif nramp = '0' and StoredData = "001011100110" then SHout <= '1' after delay1 + 742*delay_incr;
elsif nramp = '0' and StoredData = "001011100111" then SHout <= '1' after delay1 + 743*delay_incr;
elsif nramp = '0' and StoredData = "001011101000" then SHout <= '1' after delay1 + 744*delay_incr;
elsif nramp = '0' and StoredData = "001011101001" then SHout <= '1' after delay1 + 745*delay_incr;
elsif nramp = '0' and StoredData = "001011101010" then SHout <= '1' after delay1 + 746*delay_incr;
elsif nramp = '0' and StoredData = "001011101011" then SHout <= '1' after delay1 + 747*delay_incr;
elsif nramp = '0' and StoredData = "001011101100" then SHout <= '1' after delay1 + 748*delay_incr;
elsif nramp = '0' and StoredData = "001011101101" then SHout <= '1' after delay1 + 749*delay_incr;
elsif nramp = '0' and StoredData = "001011101110" then SHout <= '1' after delay1 + 750*delay_incr;
elsif nramp = '0' and StoredData = "001011101111" then SHout <= '1' after delay1 + 751*delay_incr;
elsif nramp = '0' and StoredData = "001011110000" then SHout <= '1' after delay1 + 752*delay_incr;
elsif nramp = '0' and StoredData = "001011110001" then SHout <= '1' after delay1 + 753*delay_incr;
elsif nramp = '0' and StoredData = "001011110010" then SHout <= '1' after delay1 + 754*delay_incr;
elsif nramp = '0' and StoredData = "001011110011" then SHout <= '1' after delay1 + 755*delay_incr;
elsif nramp = '0' and StoredData = "001011110100" then SHout <= '1' after delay1 + 756*delay_incr;
elsif nramp = '0' and StoredData = "001011110101" then SHout <= '1' after delay1 + 757*delay_incr;
elsif nramp = '0' and StoredData = "001011110110" then SHout <= '1' after delay1 + 758*delay_incr;
elsif nramp = '0' and StoredData = "001011110111" then SHout <= '1' after delay1 + 759*delay_incr;
elsif nramp = '0' and StoredData = "001011111000" then SHout <= '1' after delay1 + 760*delay_incr;
elsif nramp = '0' and StoredData = "001011111001" then SHout <= '1' after delay1 + 761*delay_incr;
elsif nramp = '0' and StoredData = "001011111010" then SHout <= '1' after delay1 + 762*delay_incr;
elsif nramp = '0' and StoredData = "001011111011" then SHout <= '1' after delay1 + 763*delay_incr;
elsif nramp = '0' and StoredData = "001011111100" then SHout <= '1' after delay1 + 764*delay_incr;
elsif nramp = '0' and StoredData = "001011111101" then SHout <= '1' after delay1 + 765*delay_incr;
elsif nramp = '0' and StoredData = "001011111110" then SHout <= '1' after delay1 + 766*delay_incr;
elsif nramp = '0' and StoredData = "001011111111" then SHout <= '1' after delay1 + 767*delay_incr;
elsif nramp = '0' and StoredData = "001100000000" then SHout <= '1' after delay1 + 768*delay_incr;
elsif nramp = '0' and StoredData = "001100000001" then SHout <= '1' after delay1 + 769*delay_incr;
elsif nramp = '0' and StoredData = "001100000010" then SHout <= '1' after delay1 + 770*delay_incr;
elsif nramp = '0' and StoredData = "001100000011" then SHout <= '1' after delay1 + 771*delay_incr;
elsif nramp = '0' and StoredData = "001100000100" then SHout <= '1' after delay1 + 772*delay_incr;
elsif nramp = '0' and StoredData = "001100000101" then SHout <= '1' after delay1 + 773*delay_incr;
elsif nramp = '0' and StoredData = "001100000110" then SHout <= '1' after delay1 + 774*delay_incr;
elsif nramp = '0' and StoredData = "001100000111" then SHout <= '1' after delay1 + 775*delay_incr;
elsif nramp = '0' and StoredData = "001100001000" then SHout <= '1' after delay1 + 776*delay_incr;
elsif nramp = '0' and StoredData = "001100001001" then SHout <= '1' after delay1 + 777*delay_incr;
elsif nramp = '0' and StoredData = "001100001010" then SHout <= '1' after delay1 + 778*delay_incr;
elsif nramp = '0' and StoredData = "001100001011" then SHout <= '1' after delay1 + 779*delay_incr;
elsif nramp = '0' and StoredData = "001100001100" then SHout <= '1' after delay1 + 780*delay_incr;
elsif nramp = '0' and StoredData = "001100001101" then SHout <= '1' after delay1 + 781*delay_incr;
elsif nramp = '0' and StoredData = "001100001110" then SHout <= '1' after delay1 + 782*delay_incr;
elsif nramp = '0' and StoredData = "001100001111" then SHout <= '1' after delay1 + 783*delay_incr;
elsif nramp = '0' and StoredData = "001100010000" then SHout <= '1' after delay1 + 784*delay_incr;
elsif nramp = '0' and StoredData = "001100010001" then SHout <= '1' after delay1 + 785*delay_incr;
elsif nramp = '0' and StoredData = "001100010010" then SHout <= '1' after delay1 + 786*delay_incr;
elsif nramp = '0' and StoredData = "001100010011" then SHout <= '1' after delay1 + 787*delay_incr;
elsif nramp = '0' and StoredData = "001100010100" then SHout <= '1' after delay1 + 788*delay_incr;
elsif nramp = '0' and StoredData = "001100010101" then SHout <= '1' after delay1 + 789*delay_incr;
elsif nramp = '0' and StoredData = "001100010110" then SHout <= '1' after delay1 + 790*delay_incr;
elsif nramp = '0' and StoredData = "001100010111" then SHout <= '1' after delay1 + 791*delay_incr;
elsif nramp = '0' and StoredData = "001100011000" then SHout <= '1' after delay1 + 792*delay_incr;
elsif nramp = '0' and StoredData = "001100011001" then SHout <= '1' after delay1 + 793*delay_incr;
elsif nramp = '0' and StoredData = "001100011010" then SHout <= '1' after delay1 + 794*delay_incr;
elsif nramp = '0' and StoredData = "001100011011" then SHout <= '1' after delay1 + 795*delay_incr;
elsif nramp = '0' and StoredData = "001100011100" then SHout <= '1' after delay1 + 796*delay_incr;
elsif nramp = '0' and StoredData = "001100011101" then SHout <= '1' after delay1 + 797*delay_incr;
elsif nramp = '0' and StoredData = "001100011110" then SHout <= '1' after delay1 + 798*delay_incr;
elsif nramp = '0' and StoredData = "001100011111" then SHout <= '1' after delay1 + 799*delay_incr;
elsif nramp = '0' and StoredData = "001100100000" then SHout <= '1' after delay1 + 800*delay_incr;
elsif nramp = '0' and StoredData = "001100100001" then SHout <= '1' after delay1 + 801*delay_incr;
elsif nramp = '0' and StoredData = "001100100010" then SHout <= '1' after delay1 + 802*delay_incr;
elsif nramp = '0' and StoredData = "001100100011" then SHout <= '1' after delay1 + 803*delay_incr;
elsif nramp = '0' and StoredData = "001100100100" then SHout <= '1' after delay1 + 804*delay_incr;
elsif nramp = '0' and StoredData = "001100100101" then SHout <= '1' after delay1 + 805*delay_incr;
elsif nramp = '0' and StoredData = "001100100110" then SHout <= '1' after delay1 + 806*delay_incr;
elsif nramp = '0' and StoredData = "001100100111" then SHout <= '1' after delay1 + 807*delay_incr;
elsif nramp = '0' and StoredData = "001100101000" then SHout <= '1' after delay1 + 808*delay_incr;
elsif nramp = '0' and StoredData = "001100101001" then SHout <= '1' after delay1 + 809*delay_incr;
elsif nramp = '0' and StoredData = "001100101010" then SHout <= '1' after delay1 + 810*delay_incr;
elsif nramp = '0' and StoredData = "001100101011" then SHout <= '1' after delay1 + 811*delay_incr;
elsif nramp = '0' and StoredData = "001100101100" then SHout <= '1' after delay1 + 812*delay_incr;
elsif nramp = '0' and StoredData = "001100101101" then SHout <= '1' after delay1 + 813*delay_incr;
elsif nramp = '0' and StoredData = "001100101110" then SHout <= '1' after delay1 + 814*delay_incr;
elsif nramp = '0' and StoredData = "001100101111" then SHout <= '1' after delay1 + 815*delay_incr;
elsif nramp = '0' and StoredData = "001100110000" then SHout <= '1' after delay1 + 816*delay_incr;
elsif nramp = '0' and StoredData = "001100110001" then SHout <= '1' after delay1 + 817*delay_incr;
elsif nramp = '0' and StoredData = "001100110010" then SHout <= '1' after delay1 + 818*delay_incr;
elsif nramp = '0' and StoredData = "001100110011" then SHout <= '1' after delay1 + 819*delay_incr;
elsif nramp = '0' and StoredData = "001100110100" then SHout <= '1' after delay1 + 820*delay_incr;
elsif nramp = '0' and StoredData = "001100110101" then SHout <= '1' after delay1 + 821*delay_incr;
elsif nramp = '0' and StoredData = "001100110110" then SHout <= '1' after delay1 + 822*delay_incr;
elsif nramp = '0' and StoredData = "001100110111" then SHout <= '1' after delay1 + 823*delay_incr;
elsif nramp = '0' and StoredData = "001100111000" then SHout <= '1' after delay1 + 824*delay_incr;
elsif nramp = '0' and StoredData = "001100111001" then SHout <= '1' after delay1 + 825*delay_incr;
elsif nramp = '0' and StoredData = "001100111010" then SHout <= '1' after delay1 + 826*delay_incr;
elsif nramp = '0' and StoredData = "001100111011" then SHout <= '1' after delay1 + 827*delay_incr;
elsif nramp = '0' and StoredData = "001100111100" then SHout <= '1' after delay1 + 828*delay_incr;
elsif nramp = '0' and StoredData = "001100111101" then SHout <= '1' after delay1 + 829*delay_incr;
elsif nramp = '0' and StoredData = "001100111110" then SHout <= '1' after delay1 + 830*delay_incr;
elsif nramp = '0' and StoredData = "001100111111" then SHout <= '1' after delay1 + 831*delay_incr;
elsif nramp = '0' and StoredData = "001101000000" then SHout <= '1' after delay1 + 832*delay_incr;
elsif nramp = '0' and StoredData = "001101000001" then SHout <= '1' after delay1 + 833*delay_incr;
elsif nramp = '0' and StoredData = "001101000010" then SHout <= '1' after delay1 + 834*delay_incr;
elsif nramp = '0' and StoredData = "001101000011" then SHout <= '1' after delay1 + 835*delay_incr;
elsif nramp = '0' and StoredData = "001101000100" then SHout <= '1' after delay1 + 836*delay_incr;
elsif nramp = '0' and StoredData = "001101000101" then SHout <= '1' after delay1 + 837*delay_incr;
elsif nramp = '0' and StoredData = "001101000110" then SHout <= '1' after delay1 + 838*delay_incr;
elsif nramp = '0' and StoredData = "001101000111" then SHout <= '1' after delay1 + 839*delay_incr;
elsif nramp = '0' and StoredData = "001101001000" then SHout <= '1' after delay1 + 840*delay_incr;
elsif nramp = '0' and StoredData = "001101001001" then SHout <= '1' after delay1 + 841*delay_incr;
elsif nramp = '0' and StoredData = "001101001010" then SHout <= '1' after delay1 + 842*delay_incr;
elsif nramp = '0' and StoredData = "001101001011" then SHout <= '1' after delay1 + 843*delay_incr;
elsif nramp = '0' and StoredData = "001101001100" then SHout <= '1' after delay1 + 844*delay_incr;
elsif nramp = '0' and StoredData = "001101001101" then SHout <= '1' after delay1 + 845*delay_incr;
elsif nramp = '0' and StoredData = "001101001110" then SHout <= '1' after delay1 + 846*delay_incr;
elsif nramp = '0' and StoredData = "001101001111" then SHout <= '1' after delay1 + 847*delay_incr;
elsif nramp = '0' and StoredData = "001101010000" then SHout <= '1' after delay1 + 848*delay_incr;
elsif nramp = '0' and StoredData = "001101010001" then SHout <= '1' after delay1 + 849*delay_incr;
elsif nramp = '0' and StoredData = "001101010010" then SHout <= '1' after delay1 + 850*delay_incr;
elsif nramp = '0' and StoredData = "001101010011" then SHout <= '1' after delay1 + 851*delay_incr;
elsif nramp = '0' and StoredData = "001101010100" then SHout <= '1' after delay1 + 852*delay_incr;
elsif nramp = '0' and StoredData = "001101010101" then SHout <= '1' after delay1 + 853*delay_incr;
elsif nramp = '0' and StoredData = "001101010110" then SHout <= '1' after delay1 + 854*delay_incr;
elsif nramp = '0' and StoredData = "001101010111" then SHout <= '1' after delay1 + 855*delay_incr;
elsif nramp = '0' and StoredData = "001101011000" then SHout <= '1' after delay1 + 856*delay_incr;
elsif nramp = '0' and StoredData = "001101011001" then SHout <= '1' after delay1 + 857*delay_incr;
elsif nramp = '0' and StoredData = "001101011010" then SHout <= '1' after delay1 + 858*delay_incr;
elsif nramp = '0' and StoredData = "001101011011" then SHout <= '1' after delay1 + 859*delay_incr;
elsif nramp = '0' and StoredData = "001101011100" then SHout <= '1' after delay1 + 860*delay_incr;
elsif nramp = '0' and StoredData = "001101011101" then SHout <= '1' after delay1 + 861*delay_incr;
elsif nramp = '0' and StoredData = "001101011110" then SHout <= '1' after delay1 + 862*delay_incr;
elsif nramp = '0' and StoredData = "001101011111" then SHout <= '1' after delay1 + 863*delay_incr;
elsif nramp = '0' and StoredData = "001101100000" then SHout <= '1' after delay1 + 864*delay_incr;
elsif nramp = '0' and StoredData = "001101100001" then SHout <= '1' after delay1 + 865*delay_incr;
elsif nramp = '0' and StoredData = "001101100010" then SHout <= '1' after delay1 + 866*delay_incr;
elsif nramp = '0' and StoredData = "001101100011" then SHout <= '1' after delay1 + 867*delay_incr;
elsif nramp = '0' and StoredData = "001101100100" then SHout <= '1' after delay1 + 868*delay_incr;
elsif nramp = '0' and StoredData = "001101100101" then SHout <= '1' after delay1 + 869*delay_incr;
elsif nramp = '0' and StoredData = "001101100110" then SHout <= '1' after delay1 + 870*delay_incr;
elsif nramp = '0' and StoredData = "001101100111" then SHout <= '1' after delay1 + 871*delay_incr;
elsif nramp = '0' and StoredData = "001101101000" then SHout <= '1' after delay1 + 872*delay_incr;
elsif nramp = '0' and StoredData = "001101101001" then SHout <= '1' after delay1 + 873*delay_incr;
elsif nramp = '0' and StoredData = "001101101010" then SHout <= '1' after delay1 + 874*delay_incr;
elsif nramp = '0' and StoredData = "001101101011" then SHout <= '1' after delay1 + 875*delay_incr;
elsif nramp = '0' and StoredData = "001101101100" then SHout <= '1' after delay1 + 876*delay_incr;
elsif nramp = '0' and StoredData = "001101101101" then SHout <= '1' after delay1 + 877*delay_incr;
elsif nramp = '0' and StoredData = "001101101110" then SHout <= '1' after delay1 + 878*delay_incr;
elsif nramp = '0' and StoredData = "001101101111" then SHout <= '1' after delay1 + 879*delay_incr;
elsif nramp = '0' and StoredData = "001101110000" then SHout <= '1' after delay1 + 880*delay_incr;
elsif nramp = '0' and StoredData = "001101110001" then SHout <= '1' after delay1 + 881*delay_incr;
elsif nramp = '0' and StoredData = "001101110010" then SHout <= '1' after delay1 + 882*delay_incr;
elsif nramp = '0' and StoredData = "001101110011" then SHout <= '1' after delay1 + 883*delay_incr;
elsif nramp = '0' and StoredData = "001101110100" then SHout <= '1' after delay1 + 884*delay_incr;
elsif nramp = '0' and StoredData = "001101110101" then SHout <= '1' after delay1 + 885*delay_incr;
elsif nramp = '0' and StoredData = "001101110110" then SHout <= '1' after delay1 + 886*delay_incr;
elsif nramp = '0' and StoredData = "001101110111" then SHout <= '1' after delay1 + 887*delay_incr;
elsif nramp = '0' and StoredData = "001101111000" then SHout <= '1' after delay1 + 888*delay_incr;
elsif nramp = '0' and StoredData = "001101111001" then SHout <= '1' after delay1 + 889*delay_incr;
elsif nramp = '0' and StoredData = "001101111010" then SHout <= '1' after delay1 + 890*delay_incr;
elsif nramp = '0' and StoredData = "001101111011" then SHout <= '1' after delay1 + 891*delay_incr;
elsif nramp = '0' and StoredData = "001101111100" then SHout <= '1' after delay1 + 892*delay_incr;
elsif nramp = '0' and StoredData = "001101111101" then SHout <= '1' after delay1 + 893*delay_incr;
elsif nramp = '0' and StoredData = "001101111110" then SHout <= '1' after delay1 + 894*delay_incr;
elsif nramp = '0' and StoredData = "001101111111" then SHout <= '1' after delay1 + 895*delay_incr;
elsif nramp = '0' and StoredData = "001110000000" then SHout <= '1' after delay1 + 896*delay_incr;
elsif nramp = '0' and StoredData = "001110000001" then SHout <= '1' after delay1 + 897*delay_incr;
elsif nramp = '0' and StoredData = "001110000010" then SHout <= '1' after delay1 + 898*delay_incr;
elsif nramp = '0' and StoredData = "001110000011" then SHout <= '1' after delay1 + 899*delay_incr;
elsif nramp = '0' and StoredData = "001110000100" then SHout <= '1' after delay1 + 900*delay_incr;
elsif nramp = '0' and StoredData = "001110000101" then SHout <= '1' after delay1 + 901*delay_incr;
elsif nramp = '0' and StoredData = "001110000110" then SHout <= '1' after delay1 + 902*delay_incr;
elsif nramp = '0' and StoredData = "001110000111" then SHout <= '1' after delay1 + 903*delay_incr;
elsif nramp = '0' and StoredData = "001110001000" then SHout <= '1' after delay1 + 904*delay_incr;
elsif nramp = '0' and StoredData = "001110001001" then SHout <= '1' after delay1 + 905*delay_incr;
elsif nramp = '0' and StoredData = "001110001010" then SHout <= '1' after delay1 + 906*delay_incr;
elsif nramp = '0' and StoredData = "001110001011" then SHout <= '1' after delay1 + 907*delay_incr;
elsif nramp = '0' and StoredData = "001110001100" then SHout <= '1' after delay1 + 908*delay_incr;
elsif nramp = '0' and StoredData = "001110001101" then SHout <= '1' after delay1 + 909*delay_incr;
elsif nramp = '0' and StoredData = "001110001110" then SHout <= '1' after delay1 + 910*delay_incr;
elsif nramp = '0' and StoredData = "001110001111" then SHout <= '1' after delay1 + 911*delay_incr;
elsif nramp = '0' and StoredData = "001110010000" then SHout <= '1' after delay1 + 912*delay_incr;
elsif nramp = '0' and StoredData = "001110010001" then SHout <= '1' after delay1 + 913*delay_incr;
elsif nramp = '0' and StoredData = "001110010010" then SHout <= '1' after delay1 + 914*delay_incr;
elsif nramp = '0' and StoredData = "001110010011" then SHout <= '1' after delay1 + 915*delay_incr;
elsif nramp = '0' and StoredData = "001110010100" then SHout <= '1' after delay1 + 916*delay_incr;
elsif nramp = '0' and StoredData = "001110010101" then SHout <= '1' after delay1 + 917*delay_incr;
elsif nramp = '0' and StoredData = "001110010110" then SHout <= '1' after delay1 + 918*delay_incr;
elsif nramp = '0' and StoredData = "001110010111" then SHout <= '1' after delay1 + 919*delay_incr;
elsif nramp = '0' and StoredData = "001110011000" then SHout <= '1' after delay1 + 920*delay_incr;
elsif nramp = '0' and StoredData = "001110011001" then SHout <= '1' after delay1 + 921*delay_incr;
elsif nramp = '0' and StoredData = "001110011010" then SHout <= '1' after delay1 + 922*delay_incr;
elsif nramp = '0' and StoredData = "001110011011" then SHout <= '1' after delay1 + 923*delay_incr;
elsif nramp = '0' and StoredData = "001110011100" then SHout <= '1' after delay1 + 924*delay_incr;
elsif nramp = '0' and StoredData = "001110011101" then SHout <= '1' after delay1 + 925*delay_incr;
elsif nramp = '0' and StoredData = "001110011110" then SHout <= '1' after delay1 + 926*delay_incr;
elsif nramp = '0' and StoredData = "001110011111" then SHout <= '1' after delay1 + 927*delay_incr;
elsif nramp = '0' and StoredData = "001110100000" then SHout <= '1' after delay1 + 928*delay_incr;
elsif nramp = '0' and StoredData = "001110100001" then SHout <= '1' after delay1 + 929*delay_incr;
elsif nramp = '0' and StoredData = "001110100010" then SHout <= '1' after delay1 + 930*delay_incr;
elsif nramp = '0' and StoredData = "001110100011" then SHout <= '1' after delay1 + 931*delay_incr;
elsif nramp = '0' and StoredData = "001110100100" then SHout <= '1' after delay1 + 932*delay_incr;
elsif nramp = '0' and StoredData = "001110100101" then SHout <= '1' after delay1 + 933*delay_incr;
elsif nramp = '0' and StoredData = "001110100110" then SHout <= '1' after delay1 + 934*delay_incr;
elsif nramp = '0' and StoredData = "001110100111" then SHout <= '1' after delay1 + 935*delay_incr;
elsif nramp = '0' and StoredData = "001110101000" then SHout <= '1' after delay1 + 936*delay_incr;
elsif nramp = '0' and StoredData = "001110101001" then SHout <= '1' after delay1 + 937*delay_incr;
elsif nramp = '0' and StoredData = "001110101010" then SHout <= '1' after delay1 + 938*delay_incr;
elsif nramp = '0' and StoredData = "001110101011" then SHout <= '1' after delay1 + 939*delay_incr;
elsif nramp = '0' and StoredData = "001110101100" then SHout <= '1' after delay1 + 940*delay_incr;
elsif nramp = '0' and StoredData = "001110101101" then SHout <= '1' after delay1 + 941*delay_incr;
elsif nramp = '0' and StoredData = "001110101110" then SHout <= '1' after delay1 + 942*delay_incr;
elsif nramp = '0' and StoredData = "001110101111" then SHout <= '1' after delay1 + 943*delay_incr;
elsif nramp = '0' and StoredData = "001110110000" then SHout <= '1' after delay1 + 944*delay_incr;
elsif nramp = '0' and StoredData = "001110110001" then SHout <= '1' after delay1 + 945*delay_incr;
elsif nramp = '0' and StoredData = "001110110010" then SHout <= '1' after delay1 + 946*delay_incr;
elsif nramp = '0' and StoredData = "001110110011" then SHout <= '1' after delay1 + 947*delay_incr;
elsif nramp = '0' and StoredData = "001110110100" then SHout <= '1' after delay1 + 948*delay_incr;
elsif nramp = '0' and StoredData = "001110110101" then SHout <= '1' after delay1 + 949*delay_incr;
elsif nramp = '0' and StoredData = "001110110110" then SHout <= '1' after delay1 + 950*delay_incr;
elsif nramp = '0' and StoredData = "001110110111" then SHout <= '1' after delay1 + 951*delay_incr;
elsif nramp = '0' and StoredData = "001110111000" then SHout <= '1' after delay1 + 952*delay_incr;
elsif nramp = '0' and StoredData = "001110111001" then SHout <= '1' after delay1 + 953*delay_incr;
elsif nramp = '0' and StoredData = "001110111010" then SHout <= '1' after delay1 + 954*delay_incr;
elsif nramp = '0' and StoredData = "001110111011" then SHout <= '1' after delay1 + 955*delay_incr;
elsif nramp = '0' and StoredData = "001110111100" then SHout <= '1' after delay1 + 956*delay_incr;
elsif nramp = '0' and StoredData = "001110111101" then SHout <= '1' after delay1 + 957*delay_incr;
elsif nramp = '0' and StoredData = "001110111110" then SHout <= '1' after delay1 + 958*delay_incr;
elsif nramp = '0' and StoredData = "001110111111" then SHout <= '1' after delay1 + 959*delay_incr;
elsif nramp = '0' and StoredData = "001111000000" then SHout <= '1' after delay1 + 960*delay_incr;
elsif nramp = '0' and StoredData = "001111000001" then SHout <= '1' after delay1 + 961*delay_incr;
elsif nramp = '0' and StoredData = "001111000010" then SHout <= '1' after delay1 + 962*delay_incr;
elsif nramp = '0' and StoredData = "001111000011" then SHout <= '1' after delay1 + 963*delay_incr;
elsif nramp = '0' and StoredData = "001111000100" then SHout <= '1' after delay1 + 964*delay_incr;
elsif nramp = '0' and StoredData = "001111000101" then SHout <= '1' after delay1 + 965*delay_incr;
elsif nramp = '0' and StoredData = "001111000110" then SHout <= '1' after delay1 + 966*delay_incr;
elsif nramp = '0' and StoredData = "001111000111" then SHout <= '1' after delay1 + 967*delay_incr;
elsif nramp = '0' and StoredData = "001111001000" then SHout <= '1' after delay1 + 968*delay_incr;
elsif nramp = '0' and StoredData = "001111001001" then SHout <= '1' after delay1 + 969*delay_incr;
elsif nramp = '0' and StoredData = "001111001010" then SHout <= '1' after delay1 + 970*delay_incr;
elsif nramp = '0' and StoredData = "001111001011" then SHout <= '1' after delay1 + 971*delay_incr;
elsif nramp = '0' and StoredData = "001111001100" then SHout <= '1' after delay1 + 972*delay_incr;
elsif nramp = '0' and StoredData = "001111001101" then SHout <= '1' after delay1 + 973*delay_incr;
elsif nramp = '0' and StoredData = "001111001110" then SHout <= '1' after delay1 + 974*delay_incr;
elsif nramp = '0' and StoredData = "001111001111" then SHout <= '1' after delay1 + 975*delay_incr;
elsif nramp = '0' and StoredData = "001111010000" then SHout <= '1' after delay1 + 976*delay_incr;
elsif nramp = '0' and StoredData = "001111010001" then SHout <= '1' after delay1 + 977*delay_incr;
elsif nramp = '0' and StoredData = "001111010010" then SHout <= '1' after delay1 + 978*delay_incr;
elsif nramp = '0' and StoredData = "001111010011" then SHout <= '1' after delay1 + 979*delay_incr;
elsif nramp = '0' and StoredData = "001111010100" then SHout <= '1' after delay1 + 980*delay_incr;
elsif nramp = '0' and StoredData = "001111010101" then SHout <= '1' after delay1 + 981*delay_incr;
elsif nramp = '0' and StoredData = "001111010110" then SHout <= '1' after delay1 + 982*delay_incr;
elsif nramp = '0' and StoredData = "001111010111" then SHout <= '1' after delay1 + 983*delay_incr;
elsif nramp = '0' and StoredData = "001111011000" then SHout <= '1' after delay1 + 984*delay_incr;
elsif nramp = '0' and StoredData = "001111011001" then SHout <= '1' after delay1 + 985*delay_incr;
elsif nramp = '0' and StoredData = "001111011010" then SHout <= '1' after delay1 + 986*delay_incr;
elsif nramp = '0' and StoredData = "001111011011" then SHout <= '1' after delay1 + 987*delay_incr;
elsif nramp = '0' and StoredData = "001111011100" then SHout <= '1' after delay1 + 988*delay_incr;
elsif nramp = '0' and StoredData = "001111011101" then SHout <= '1' after delay1 + 989*delay_incr;
elsif nramp = '0' and StoredData = "001111011110" then SHout <= '1' after delay1 + 990*delay_incr;
elsif nramp = '0' and StoredData = "001111011111" then SHout <= '1' after delay1 + 991*delay_incr;
elsif nramp = '0' and StoredData = "001111100000" then SHout <= '1' after delay1 + 992*delay_incr;
elsif nramp = '0' and StoredData = "001111100001" then SHout <= '1' after delay1 + 993*delay_incr;
elsif nramp = '0' and StoredData = "001111100010" then SHout <= '1' after delay1 + 994*delay_incr;
elsif nramp = '0' and StoredData = "001111100011" then SHout <= '1' after delay1 + 995*delay_incr;
elsif nramp = '0' and StoredData = "001111100100" then SHout <= '1' after delay1 + 996*delay_incr;
elsif nramp = '0' and StoredData = "001111100101" then SHout <= '1' after delay1 + 997*delay_incr;
elsif nramp = '0' and StoredData = "001111100110" then SHout <= '1' after delay1 + 998*delay_incr;
elsif nramp = '0' and StoredData = "001111100111" then SHout <= '1' after delay1 + 999*delay_incr;
elsif nramp = '0' and StoredData = "001111101000" then SHout <= '1' after delay1 + 1000*delay_incr;
elsif nramp = '0' and StoredData = "001111101001" then SHout <= '1' after delay1 + 1001*delay_incr;
elsif nramp = '0' and StoredData = "001111101010" then SHout <= '1' after delay1 + 1002*delay_incr;
elsif nramp = '0' and StoredData = "001111101011" then SHout <= '1' after delay1 + 1003*delay_incr;
elsif nramp = '0' and StoredData = "001111101100" then SHout <= '1' after delay1 + 1004*delay_incr;
elsif nramp = '0' and StoredData = "001111101101" then SHout <= '1' after delay1 + 1005*delay_incr;
elsif nramp = '0' and StoredData = "001111101110" then SHout <= '1' after delay1 + 1006*delay_incr;
elsif nramp = '0' and StoredData = "001111101111" then SHout <= '1' after delay1 + 1007*delay_incr;
elsif nramp = '0' and StoredData = "001111110000" then SHout <= '1' after delay1 + 1008*delay_incr;
elsif nramp = '0' and StoredData = "001111110001" then SHout <= '1' after delay1 + 1009*delay_incr;
elsif nramp = '0' and StoredData = "001111110010" then SHout <= '1' after delay1 + 1010*delay_incr;
elsif nramp = '0' and StoredData = "001111110011" then SHout <= '1' after delay1 + 1011*delay_incr;
elsif nramp = '0' and StoredData = "001111110100" then SHout <= '1' after delay1 + 1012*delay_incr;
elsif nramp = '0' and StoredData = "001111110101" then SHout <= '1' after delay1 + 1013*delay_incr;
elsif nramp = '0' and StoredData = "001111110110" then SHout <= '1' after delay1 + 1014*delay_incr;
elsif nramp = '0' and StoredData = "001111110111" then SHout <= '1' after delay1 + 1015*delay_incr;
elsif nramp = '0' and StoredData = "001111111000" then SHout <= '1' after delay1 + 1016*delay_incr;
elsif nramp = '0' and StoredData = "001111111001" then SHout <= '1' after delay1 + 1017*delay_incr;
elsif nramp = '0' and StoredData = "001111111010" then SHout <= '1' after delay1 + 1018*delay_incr;
elsif nramp = '0' and StoredData = "001111111011" then SHout <= '1' after delay1 + 1019*delay_incr;
elsif nramp = '0' and StoredData = "001111111100" then SHout <= '1' after delay1 + 1020*delay_incr;
elsif nramp = '0' and StoredData = "001111111101" then SHout <= '1' after delay1 + 1021*delay_incr;
elsif nramp = '0' and StoredData = "001111111110" then SHout <= '1' after delay1 + 1022*delay_incr;
elsif nramp = '0' and StoredData = "001111111111" then SHout <= '1' after delay1 + 1023*delay_incr;
elsif nramp = '0' and StoredData = "010000000000" then SHout <= '1' after delay1 + 1024*delay_incr;
elsif nramp = '0' and StoredData = "010000000001" then SHout <= '1' after delay1 + 1025*delay_incr;
elsif nramp = '0' and StoredData = "010000000010" then SHout <= '1' after delay1 + 1026*delay_incr;
elsif nramp = '0' and StoredData = "010000000011" then SHout <= '1' after delay1 + 1027*delay_incr;
elsif nramp = '0' and StoredData = "010000000100" then SHout <= '1' after delay1 + 1028*delay_incr;
elsif nramp = '0' and StoredData = "010000000101" then SHout <= '1' after delay1 + 1029*delay_incr;
elsif nramp = '0' and StoredData = "010000000110" then SHout <= '1' after delay1 + 1030*delay_incr;
elsif nramp = '0' and StoredData = "010000000111" then SHout <= '1' after delay1 + 1031*delay_incr;
elsif nramp = '0' and StoredData = "010000001000" then SHout <= '1' after delay1 + 1032*delay_incr;
elsif nramp = '0' and StoredData = "010000001001" then SHout <= '1' after delay1 + 1033*delay_incr;
elsif nramp = '0' and StoredData = "010000001010" then SHout <= '1' after delay1 + 1034*delay_incr;
elsif nramp = '0' and StoredData = "010000001011" then SHout <= '1' after delay1 + 1035*delay_incr;
elsif nramp = '0' and StoredData = "010000001100" then SHout <= '1' after delay1 + 1036*delay_incr;
elsif nramp = '0' and StoredData = "010000001101" then SHout <= '1' after delay1 + 1037*delay_incr;
elsif nramp = '0' and StoredData = "010000001110" then SHout <= '1' after delay1 + 1038*delay_incr;
elsif nramp = '0' and StoredData = "010000001111" then SHout <= '1' after delay1 + 1039*delay_incr;
elsif nramp = '0' and StoredData = "010000010000" then SHout <= '1' after delay1 + 1040*delay_incr;
elsif nramp = '0' and StoredData = "010000010001" then SHout <= '1' after delay1 + 1041*delay_incr;
elsif nramp = '0' and StoredData = "010000010010" then SHout <= '1' after delay1 + 1042*delay_incr;
elsif nramp = '0' and StoredData = "010000010011" then SHout <= '1' after delay1 + 1043*delay_incr;
elsif nramp = '0' and StoredData = "010000010100" then SHout <= '1' after delay1 + 1044*delay_incr;
elsif nramp = '0' and StoredData = "010000010101" then SHout <= '1' after delay1 + 1045*delay_incr;
elsif nramp = '0' and StoredData = "010000010110" then SHout <= '1' after delay1 + 1046*delay_incr;
elsif nramp = '0' and StoredData = "010000010111" then SHout <= '1' after delay1 + 1047*delay_incr;
elsif nramp = '0' and StoredData = "010000011000" then SHout <= '1' after delay1 + 1048*delay_incr;
elsif nramp = '0' and StoredData = "010000011001" then SHout <= '1' after delay1 + 1049*delay_incr;
elsif nramp = '0' and StoredData = "010000011010" then SHout <= '1' after delay1 + 1050*delay_incr;
elsif nramp = '0' and StoredData = "010000011011" then SHout <= '1' after delay1 + 1051*delay_incr;
elsif nramp = '0' and StoredData = "010000011100" then SHout <= '1' after delay1 + 1052*delay_incr;
elsif nramp = '0' and StoredData = "010000011101" then SHout <= '1' after delay1 + 1053*delay_incr;
elsif nramp = '0' and StoredData = "010000011110" then SHout <= '1' after delay1 + 1054*delay_incr;
elsif nramp = '0' and StoredData = "010000011111" then SHout <= '1' after delay1 + 1055*delay_incr;
elsif nramp = '0' and StoredData = "010000100000" then SHout <= '1' after delay1 + 1056*delay_incr;
elsif nramp = '0' and StoredData = "010000100001" then SHout <= '1' after delay1 + 1057*delay_incr;
elsif nramp = '0' and StoredData = "010000100010" then SHout <= '1' after delay1 + 1058*delay_incr;
elsif nramp = '0' and StoredData = "010000100011" then SHout <= '1' after delay1 + 1059*delay_incr;
elsif nramp = '0' and StoredData = "010000100100" then SHout <= '1' after delay1 + 1060*delay_incr;
elsif nramp = '0' and StoredData = "010000100101" then SHout <= '1' after delay1 + 1061*delay_incr;
elsif nramp = '0' and StoredData = "010000100110" then SHout <= '1' after delay1 + 1062*delay_incr;
elsif nramp = '0' and StoredData = "010000100111" then SHout <= '1' after delay1 + 1063*delay_incr;
elsif nramp = '0' and StoredData = "010000101000" then SHout <= '1' after delay1 + 1064*delay_incr;
elsif nramp = '0' and StoredData = "010000101001" then SHout <= '1' after delay1 + 1065*delay_incr;
elsif nramp = '0' and StoredData = "010000101010" then SHout <= '1' after delay1 + 1066*delay_incr;
elsif nramp = '0' and StoredData = "010000101011" then SHout <= '1' after delay1 + 1067*delay_incr;
elsif nramp = '0' and StoredData = "010000101100" then SHout <= '1' after delay1 + 1068*delay_incr;
elsif nramp = '0' and StoredData = "010000101101" then SHout <= '1' after delay1 + 1069*delay_incr;
elsif nramp = '0' and StoredData = "010000101110" then SHout <= '1' after delay1 + 1070*delay_incr;
elsif nramp = '0' and StoredData = "010000101111" then SHout <= '1' after delay1 + 1071*delay_incr;
elsif nramp = '0' and StoredData = "010000110000" then SHout <= '1' after delay1 + 1072*delay_incr;
elsif nramp = '0' and StoredData = "010000110001" then SHout <= '1' after delay1 + 1073*delay_incr;
elsif nramp = '0' and StoredData = "010000110010" then SHout <= '1' after delay1 + 1074*delay_incr;
elsif nramp = '0' and StoredData = "010000110011" then SHout <= '1' after delay1 + 1075*delay_incr;
elsif nramp = '0' and StoredData = "010000110100" then SHout <= '1' after delay1 + 1076*delay_incr;
elsif nramp = '0' and StoredData = "010000110101" then SHout <= '1' after delay1 + 1077*delay_incr;
elsif nramp = '0' and StoredData = "010000110110" then SHout <= '1' after delay1 + 1078*delay_incr;
elsif nramp = '0' and StoredData = "010000110111" then SHout <= '1' after delay1 + 1079*delay_incr;
elsif nramp = '0' and StoredData = "010000111000" then SHout <= '1' after delay1 + 1080*delay_incr;
elsif nramp = '0' and StoredData = "010000111001" then SHout <= '1' after delay1 + 1081*delay_incr;
elsif nramp = '0' and StoredData = "010000111010" then SHout <= '1' after delay1 + 1082*delay_incr;
elsif nramp = '0' and StoredData = "010000111011" then SHout <= '1' after delay1 + 1083*delay_incr;
elsif nramp = '0' and StoredData = "010000111100" then SHout <= '1' after delay1 + 1084*delay_incr;
elsif nramp = '0' and StoredData = "010000111101" then SHout <= '1' after delay1 + 1085*delay_incr;
elsif nramp = '0' and StoredData = "010000111110" then SHout <= '1' after delay1 + 1086*delay_incr;
elsif nramp = '0' and StoredData = "010000111111" then SHout <= '1' after delay1 + 1087*delay_incr;
elsif nramp = '0' and StoredData = "010001000000" then SHout <= '1' after delay1 + 1088*delay_incr;
elsif nramp = '0' and StoredData = "010001000001" then SHout <= '1' after delay1 + 1089*delay_incr;
elsif nramp = '0' and StoredData = "010001000010" then SHout <= '1' after delay1 + 1090*delay_incr;
elsif nramp = '0' and StoredData = "010001000011" then SHout <= '1' after delay1 + 1091*delay_incr;
elsif nramp = '0' and StoredData = "010001000100" then SHout <= '1' after delay1 + 1092*delay_incr;
elsif nramp = '0' and StoredData = "010001000101" then SHout <= '1' after delay1 + 1093*delay_incr;
elsif nramp = '0' and StoredData = "010001000110" then SHout <= '1' after delay1 + 1094*delay_incr;
elsif nramp = '0' and StoredData = "010001000111" then SHout <= '1' after delay1 + 1095*delay_incr;
elsif nramp = '0' and StoredData = "010001001000" then SHout <= '1' after delay1 + 1096*delay_incr;
elsif nramp = '0' and StoredData = "010001001001" then SHout <= '1' after delay1 + 1097*delay_incr;
elsif nramp = '0' and StoredData = "010001001010" then SHout <= '1' after delay1 + 1098*delay_incr;
elsif nramp = '0' and StoredData = "010001001011" then SHout <= '1' after delay1 + 1099*delay_incr;
elsif nramp = '0' and StoredData = "010001001100" then SHout <= '1' after delay1 + 1100*delay_incr;
elsif nramp = '0' and StoredData = "010001001101" then SHout <= '1' after delay1 + 1101*delay_incr;
elsif nramp = '0' and StoredData = "010001001110" then SHout <= '1' after delay1 + 1102*delay_incr;
elsif nramp = '0' and StoredData = "010001001111" then SHout <= '1' after delay1 + 1103*delay_incr;
elsif nramp = '0' and StoredData = "010001010000" then SHout <= '1' after delay1 + 1104*delay_incr;
elsif nramp = '0' and StoredData = "010001010001" then SHout <= '1' after delay1 + 1105*delay_incr;
elsif nramp = '0' and StoredData = "010001010010" then SHout <= '1' after delay1 + 1106*delay_incr;
elsif nramp = '0' and StoredData = "010001010011" then SHout <= '1' after delay1 + 1107*delay_incr;
elsif nramp = '0' and StoredData = "010001010100" then SHout <= '1' after delay1 + 1108*delay_incr;
elsif nramp = '0' and StoredData = "010001010101" then SHout <= '1' after delay1 + 1109*delay_incr;
elsif nramp = '0' and StoredData = "010001010110" then SHout <= '1' after delay1 + 1110*delay_incr;
elsif nramp = '0' and StoredData = "010001010111" then SHout <= '1' after delay1 + 1111*delay_incr;
elsif nramp = '0' and StoredData = "010001011000" then SHout <= '1' after delay1 + 1112*delay_incr;
elsif nramp = '0' and StoredData = "010001011001" then SHout <= '1' after delay1 + 1113*delay_incr;
elsif nramp = '0' and StoredData = "010001011010" then SHout <= '1' after delay1 + 1114*delay_incr;
elsif nramp = '0' and StoredData = "010001011011" then SHout <= '1' after delay1 + 1115*delay_incr;
elsif nramp = '0' and StoredData = "010001011100" then SHout <= '1' after delay1 + 1116*delay_incr;
elsif nramp = '0' and StoredData = "010001011101" then SHout <= '1' after delay1 + 1117*delay_incr;
elsif nramp = '0' and StoredData = "010001011110" then SHout <= '1' after delay1 + 1118*delay_incr;
elsif nramp = '0' and StoredData = "010001011111" then SHout <= '1' after delay1 + 1119*delay_incr;
elsif nramp = '0' and StoredData = "010001100000" then SHout <= '1' after delay1 + 1120*delay_incr;
elsif nramp = '0' and StoredData = "010001100001" then SHout <= '1' after delay1 + 1121*delay_incr;
elsif nramp = '0' and StoredData = "010001100010" then SHout <= '1' after delay1 + 1122*delay_incr;
elsif nramp = '0' and StoredData = "010001100011" then SHout <= '1' after delay1 + 1123*delay_incr;
elsif nramp = '0' and StoredData = "010001100100" then SHout <= '1' after delay1 + 1124*delay_incr;
elsif nramp = '0' and StoredData = "010001100101" then SHout <= '1' after delay1 + 1125*delay_incr;
elsif nramp = '0' and StoredData = "010001100110" then SHout <= '1' after delay1 + 1126*delay_incr;
elsif nramp = '0' and StoredData = "010001100111" then SHout <= '1' after delay1 + 1127*delay_incr;
elsif nramp = '0' and StoredData = "010001101000" then SHout <= '1' after delay1 + 1128*delay_incr;
elsif nramp = '0' and StoredData = "010001101001" then SHout <= '1' after delay1 + 1129*delay_incr;
elsif nramp = '0' and StoredData = "010001101010" then SHout <= '1' after delay1 + 1130*delay_incr;
elsif nramp = '0' and StoredData = "010001101011" then SHout <= '1' after delay1 + 1131*delay_incr;
elsif nramp = '0' and StoredData = "010001101100" then SHout <= '1' after delay1 + 1132*delay_incr;
elsif nramp = '0' and StoredData = "010001101101" then SHout <= '1' after delay1 + 1133*delay_incr;
elsif nramp = '0' and StoredData = "010001101110" then SHout <= '1' after delay1 + 1134*delay_incr;
elsif nramp = '0' and StoredData = "010001101111" then SHout <= '1' after delay1 + 1135*delay_incr;
elsif nramp = '0' and StoredData = "010001110000" then SHout <= '1' after delay1 + 1136*delay_incr;
elsif nramp = '0' and StoredData = "010001110001" then SHout <= '1' after delay1 + 1137*delay_incr;
elsif nramp = '0' and StoredData = "010001110010" then SHout <= '1' after delay1 + 1138*delay_incr;
elsif nramp = '0' and StoredData = "010001110011" then SHout <= '1' after delay1 + 1139*delay_incr;
elsif nramp = '0' and StoredData = "010001110100" then SHout <= '1' after delay1 + 1140*delay_incr;
elsif nramp = '0' and StoredData = "010001110101" then SHout <= '1' after delay1 + 1141*delay_incr;
elsif nramp = '0' and StoredData = "010001110110" then SHout <= '1' after delay1 + 1142*delay_incr;
elsif nramp = '0' and StoredData = "010001110111" then SHout <= '1' after delay1 + 1143*delay_incr;
elsif nramp = '0' and StoredData = "010001111000" then SHout <= '1' after delay1 + 1144*delay_incr;
elsif nramp = '0' and StoredData = "010001111001" then SHout <= '1' after delay1 + 1145*delay_incr;
elsif nramp = '0' and StoredData = "010001111010" then SHout <= '1' after delay1 + 1146*delay_incr;
elsif nramp = '0' and StoredData = "010001111011" then SHout <= '1' after delay1 + 1147*delay_incr;
elsif nramp = '0' and StoredData = "010001111100" then SHout <= '1' after delay1 + 1148*delay_incr;
elsif nramp = '0' and StoredData = "010001111101" then SHout <= '1' after delay1 + 1149*delay_incr;
elsif nramp = '0' and StoredData = "010001111110" then SHout <= '1' after delay1 + 1150*delay_incr;
elsif nramp = '0' and StoredData = "010001111111" then SHout <= '1' after delay1 + 1151*delay_incr;
elsif nramp = '0' and StoredData = "010010000000" then SHout <= '1' after delay1 + 1152*delay_incr;
elsif nramp = '0' and StoredData = "010010000001" then SHout <= '1' after delay1 + 1153*delay_incr;
elsif nramp = '0' and StoredData = "010010000010" then SHout <= '1' after delay1 + 1154*delay_incr;
elsif nramp = '0' and StoredData = "010010000011" then SHout <= '1' after delay1 + 1155*delay_incr;
elsif nramp = '0' and StoredData = "010010000100" then SHout <= '1' after delay1 + 1156*delay_incr;
elsif nramp = '0' and StoredData = "010010000101" then SHout <= '1' after delay1 + 1157*delay_incr;
elsif nramp = '0' and StoredData = "010010000110" then SHout <= '1' after delay1 + 1158*delay_incr;
elsif nramp = '0' and StoredData = "010010000111" then SHout <= '1' after delay1 + 1159*delay_incr;
elsif nramp = '0' and StoredData = "010010001000" then SHout <= '1' after delay1 + 1160*delay_incr;
elsif nramp = '0' and StoredData = "010010001001" then SHout <= '1' after delay1 + 1161*delay_incr;
elsif nramp = '0' and StoredData = "010010001010" then SHout <= '1' after delay1 + 1162*delay_incr;
elsif nramp = '0' and StoredData = "010010001011" then SHout <= '1' after delay1 + 1163*delay_incr;
elsif nramp = '0' and StoredData = "010010001100" then SHout <= '1' after delay1 + 1164*delay_incr;
elsif nramp = '0' and StoredData = "010010001101" then SHout <= '1' after delay1 + 1165*delay_incr;
elsif nramp = '0' and StoredData = "010010001110" then SHout <= '1' after delay1 + 1166*delay_incr;
elsif nramp = '0' and StoredData = "010010001111" then SHout <= '1' after delay1 + 1167*delay_incr;
elsif nramp = '0' and StoredData = "010010010000" then SHout <= '1' after delay1 + 1168*delay_incr;
elsif nramp = '0' and StoredData = "010010010001" then SHout <= '1' after delay1 + 1169*delay_incr;
elsif nramp = '0' and StoredData = "010010010010" then SHout <= '1' after delay1 + 1170*delay_incr;
elsif nramp = '0' and StoredData = "010010010011" then SHout <= '1' after delay1 + 1171*delay_incr;
elsif nramp = '0' and StoredData = "010010010100" then SHout <= '1' after delay1 + 1172*delay_incr;
elsif nramp = '0' and StoredData = "010010010101" then SHout <= '1' after delay1 + 1173*delay_incr;
elsif nramp = '0' and StoredData = "010010010110" then SHout <= '1' after delay1 + 1174*delay_incr;
elsif nramp = '0' and StoredData = "010010010111" then SHout <= '1' after delay1 + 1175*delay_incr;
elsif nramp = '0' and StoredData = "010010011000" then SHout <= '1' after delay1 + 1176*delay_incr;
elsif nramp = '0' and StoredData = "010010011001" then SHout <= '1' after delay1 + 1177*delay_incr;
elsif nramp = '0' and StoredData = "010010011010" then SHout <= '1' after delay1 + 1178*delay_incr;
elsif nramp = '0' and StoredData = "010010011011" then SHout <= '1' after delay1 + 1179*delay_incr;
elsif nramp = '0' and StoredData = "010010011100" then SHout <= '1' after delay1 + 1180*delay_incr;
elsif nramp = '0' and StoredData = "010010011101" then SHout <= '1' after delay1 + 1181*delay_incr;
elsif nramp = '0' and StoredData = "010010011110" then SHout <= '1' after delay1 + 1182*delay_incr;
elsif nramp = '0' and StoredData = "010010011111" then SHout <= '1' after delay1 + 1183*delay_incr;
elsif nramp = '0' and StoredData = "010010100000" then SHout <= '1' after delay1 + 1184*delay_incr;
elsif nramp = '0' and StoredData = "010010100001" then SHout <= '1' after delay1 + 1185*delay_incr;
elsif nramp = '0' and StoredData = "010010100010" then SHout <= '1' after delay1 + 1186*delay_incr;
elsif nramp = '0' and StoredData = "010010100011" then SHout <= '1' after delay1 + 1187*delay_incr;
elsif nramp = '0' and StoredData = "010010100100" then SHout <= '1' after delay1 + 1188*delay_incr;
elsif nramp = '0' and StoredData = "010010100101" then SHout <= '1' after delay1 + 1189*delay_incr;
elsif nramp = '0' and StoredData = "010010100110" then SHout <= '1' after delay1 + 1190*delay_incr;
elsif nramp = '0' and StoredData = "010010100111" then SHout <= '1' after delay1 + 1191*delay_incr;
elsif nramp = '0' and StoredData = "010010101000" then SHout <= '1' after delay1 + 1192*delay_incr;
elsif nramp = '0' and StoredData = "010010101001" then SHout <= '1' after delay1 + 1193*delay_incr;
elsif nramp = '0' and StoredData = "010010101010" then SHout <= '1' after delay1 + 1194*delay_incr;
elsif nramp = '0' and StoredData = "010010101011" then SHout <= '1' after delay1 + 1195*delay_incr;
elsif nramp = '0' and StoredData = "010010101100" then SHout <= '1' after delay1 + 1196*delay_incr;
elsif nramp = '0' and StoredData = "010010101101" then SHout <= '1' after delay1 + 1197*delay_incr;
elsif nramp = '0' and StoredData = "010010101110" then SHout <= '1' after delay1 + 1198*delay_incr;
elsif nramp = '0' and StoredData = "010010101111" then SHout <= '1' after delay1 + 1199*delay_incr;
elsif nramp = '0' and StoredData = "010010110000" then SHout <= '1' after delay1 + 1200*delay_incr;
elsif nramp = '0' and StoredData = "010010110001" then SHout <= '1' after delay1 + 1201*delay_incr;
elsif nramp = '0' and StoredData = "010010110010" then SHout <= '1' after delay1 + 1202*delay_incr;
elsif nramp = '0' and StoredData = "010010110011" then SHout <= '1' after delay1 + 1203*delay_incr;
elsif nramp = '0' and StoredData = "010010110100" then SHout <= '1' after delay1 + 1204*delay_incr;
elsif nramp = '0' and StoredData = "010010110101" then SHout <= '1' after delay1 + 1205*delay_incr;
elsif nramp = '0' and StoredData = "010010110110" then SHout <= '1' after delay1 + 1206*delay_incr;
elsif nramp = '0' and StoredData = "010010110111" then SHout <= '1' after delay1 + 1207*delay_incr;
elsif nramp = '0' and StoredData = "010010111000" then SHout <= '1' after delay1 + 1208*delay_incr;
elsif nramp = '0' and StoredData = "010010111001" then SHout <= '1' after delay1 + 1209*delay_incr;
elsif nramp = '0' and StoredData = "010010111010" then SHout <= '1' after delay1 + 1210*delay_incr;
elsif nramp = '0' and StoredData = "010010111011" then SHout <= '1' after delay1 + 1211*delay_incr;
elsif nramp = '0' and StoredData = "010010111100" then SHout <= '1' after delay1 + 1212*delay_incr;
elsif nramp = '0' and StoredData = "010010111101" then SHout <= '1' after delay1 + 1213*delay_incr;
elsif nramp = '0' and StoredData = "010010111110" then SHout <= '1' after delay1 + 1214*delay_incr;
elsif nramp = '0' and StoredData = "010010111111" then SHout <= '1' after delay1 + 1215*delay_incr;
elsif nramp = '0' and StoredData = "010011000000" then SHout <= '1' after delay1 + 1216*delay_incr;
elsif nramp = '0' and StoredData = "010011000001" then SHout <= '1' after delay1 + 1217*delay_incr;
elsif nramp = '0' and StoredData = "010011000010" then SHout <= '1' after delay1 + 1218*delay_incr;
elsif nramp = '0' and StoredData = "010011000011" then SHout <= '1' after delay1 + 1219*delay_incr;
elsif nramp = '0' and StoredData = "010011000100" then SHout <= '1' after delay1 + 1220*delay_incr;
elsif nramp = '0' and StoredData = "010011000101" then SHout <= '1' after delay1 + 1221*delay_incr;
elsif nramp = '0' and StoredData = "010011000110" then SHout <= '1' after delay1 + 1222*delay_incr;
elsif nramp = '0' and StoredData = "010011000111" then SHout <= '1' after delay1 + 1223*delay_incr;
elsif nramp = '0' and StoredData = "010011001000" then SHout <= '1' after delay1 + 1224*delay_incr;
elsif nramp = '0' and StoredData = "010011001001" then SHout <= '1' after delay1 + 1225*delay_incr;
elsif nramp = '0' and StoredData = "010011001010" then SHout <= '1' after delay1 + 1226*delay_incr;
elsif nramp = '0' and StoredData = "010011001011" then SHout <= '1' after delay1 + 1227*delay_incr;
elsif nramp = '0' and StoredData = "010011001100" then SHout <= '1' after delay1 + 1228*delay_incr;
elsif nramp = '0' and StoredData = "010011001101" then SHout <= '1' after delay1 + 1229*delay_incr;
elsif nramp = '0' and StoredData = "010011001110" then SHout <= '1' after delay1 + 1230*delay_incr;
elsif nramp = '0' and StoredData = "010011001111" then SHout <= '1' after delay1 + 1231*delay_incr;
elsif nramp = '0' and StoredData = "010011010000" then SHout <= '1' after delay1 + 1232*delay_incr;
elsif nramp = '0' and StoredData = "010011010001" then SHout <= '1' after delay1 + 1233*delay_incr;
elsif nramp = '0' and StoredData = "010011010010" then SHout <= '1' after delay1 + 1234*delay_incr;
elsif nramp = '0' and StoredData = "010011010011" then SHout <= '1' after delay1 + 1235*delay_incr;
elsif nramp = '0' and StoredData = "010011010100" then SHout <= '1' after delay1 + 1236*delay_incr;
elsif nramp = '0' and StoredData = "010011010101" then SHout <= '1' after delay1 + 1237*delay_incr;
elsif nramp = '0' and StoredData = "010011010110" then SHout <= '1' after delay1 + 1238*delay_incr;
elsif nramp = '0' and StoredData = "010011010111" then SHout <= '1' after delay1 + 1239*delay_incr;
elsif nramp = '0' and StoredData = "010011011000" then SHout <= '1' after delay1 + 1240*delay_incr;
elsif nramp = '0' and StoredData = "010011011001" then SHout <= '1' after delay1 + 1241*delay_incr;
elsif nramp = '0' and StoredData = "010011011010" then SHout <= '1' after delay1 + 1242*delay_incr;
elsif nramp = '0' and StoredData = "010011011011" then SHout <= '1' after delay1 + 1243*delay_incr;
elsif nramp = '0' and StoredData = "010011011100" then SHout <= '1' after delay1 + 1244*delay_incr;
elsif nramp = '0' and StoredData = "010011011101" then SHout <= '1' after delay1 + 1245*delay_incr;
elsif nramp = '0' and StoredData = "010011011110" then SHout <= '1' after delay1 + 1246*delay_incr;
elsif nramp = '0' and StoredData = "010011011111" then SHout <= '1' after delay1 + 1247*delay_incr;
elsif nramp = '0' and StoredData = "010011100000" then SHout <= '1' after delay1 + 1248*delay_incr;
elsif nramp = '0' and StoredData = "010011100001" then SHout <= '1' after delay1 + 1249*delay_incr;
elsif nramp = '0' and StoredData = "010011100010" then SHout <= '1' after delay1 + 1250*delay_incr;
elsif nramp = '0' and StoredData = "010011100011" then SHout <= '1' after delay1 + 1251*delay_incr;
elsif nramp = '0' and StoredData = "010011100100" then SHout <= '1' after delay1 + 1252*delay_incr;
elsif nramp = '0' and StoredData = "010011100101" then SHout <= '1' after delay1 + 1253*delay_incr;
elsif nramp = '0' and StoredData = "010011100110" then SHout <= '1' after delay1 + 1254*delay_incr;
elsif nramp = '0' and StoredData = "010011100111" then SHout <= '1' after delay1 + 1255*delay_incr;
elsif nramp = '0' and StoredData = "010011101000" then SHout <= '1' after delay1 + 1256*delay_incr;
elsif nramp = '0' and StoredData = "010011101001" then SHout <= '1' after delay1 + 1257*delay_incr;
elsif nramp = '0' and StoredData = "010011101010" then SHout <= '1' after delay1 + 1258*delay_incr;
elsif nramp = '0' and StoredData = "010011101011" then SHout <= '1' after delay1 + 1259*delay_incr;
elsif nramp = '0' and StoredData = "010011101100" then SHout <= '1' after delay1 + 1260*delay_incr;
elsif nramp = '0' and StoredData = "010011101101" then SHout <= '1' after delay1 + 1261*delay_incr;
elsif nramp = '0' and StoredData = "010011101110" then SHout <= '1' after delay1 + 1262*delay_incr;
elsif nramp = '0' and StoredData = "010011101111" then SHout <= '1' after delay1 + 1263*delay_incr;
elsif nramp = '0' and StoredData = "010011110000" then SHout <= '1' after delay1 + 1264*delay_incr;
elsif nramp = '0' and StoredData = "010011110001" then SHout <= '1' after delay1 + 1265*delay_incr;
elsif nramp = '0' and StoredData = "010011110010" then SHout <= '1' after delay1 + 1266*delay_incr;
elsif nramp = '0' and StoredData = "010011110011" then SHout <= '1' after delay1 + 1267*delay_incr;
elsif nramp = '0' and StoredData = "010011110100" then SHout <= '1' after delay1 + 1268*delay_incr;
elsif nramp = '0' and StoredData = "010011110101" then SHout <= '1' after delay1 + 1269*delay_incr;
elsif nramp = '0' and StoredData = "010011110110" then SHout <= '1' after delay1 + 1270*delay_incr;
elsif nramp = '0' and StoredData = "010011110111" then SHout <= '1' after delay1 + 1271*delay_incr;
elsif nramp = '0' and StoredData = "010011111000" then SHout <= '1' after delay1 + 1272*delay_incr;
elsif nramp = '0' and StoredData = "010011111001" then SHout <= '1' after delay1 + 1273*delay_incr;
elsif nramp = '0' and StoredData = "010011111010" then SHout <= '1' after delay1 + 1274*delay_incr;
elsif nramp = '0' and StoredData = "010011111011" then SHout <= '1' after delay1 + 1275*delay_incr;
elsif nramp = '0' and StoredData = "010011111100" then SHout <= '1' after delay1 + 1276*delay_incr;
elsif nramp = '0' and StoredData = "010011111101" then SHout <= '1' after delay1 + 1277*delay_incr;
elsif nramp = '0' and StoredData = "010011111110" then SHout <= '1' after delay1 + 1278*delay_incr;
elsif nramp = '0' and StoredData = "010011111111" then SHout <= '1' after delay1 + 1279*delay_incr;
elsif nramp = '0' and StoredData = "010100000000" then SHout <= '1' after delay1 + 1280*delay_incr;
elsif nramp = '0' and StoredData = "010100000001" then SHout <= '1' after delay1 + 1281*delay_incr;
elsif nramp = '0' and StoredData = "010100000010" then SHout <= '1' after delay1 + 1282*delay_incr;
elsif nramp = '0' and StoredData = "010100000011" then SHout <= '1' after delay1 + 1283*delay_incr;
elsif nramp = '0' and StoredData = "010100000100" then SHout <= '1' after delay1 + 1284*delay_incr;
elsif nramp = '0' and StoredData = "010100000101" then SHout <= '1' after delay1 + 1285*delay_incr;
elsif nramp = '0' and StoredData = "010100000110" then SHout <= '1' after delay1 + 1286*delay_incr;
elsif nramp = '0' and StoredData = "010100000111" then SHout <= '1' after delay1 + 1287*delay_incr;
elsif nramp = '0' and StoredData = "010100001000" then SHout <= '1' after delay1 + 1288*delay_incr;
elsif nramp = '0' and StoredData = "010100001001" then SHout <= '1' after delay1 + 1289*delay_incr;
elsif nramp = '0' and StoredData = "010100001010" then SHout <= '1' after delay1 + 1290*delay_incr;
elsif nramp = '0' and StoredData = "010100001011" then SHout <= '1' after delay1 + 1291*delay_incr;
elsif nramp = '0' and StoredData = "010100001100" then SHout <= '1' after delay1 + 1292*delay_incr;
elsif nramp = '0' and StoredData = "010100001101" then SHout <= '1' after delay1 + 1293*delay_incr;
elsif nramp = '0' and StoredData = "010100001110" then SHout <= '1' after delay1 + 1294*delay_incr;
elsif nramp = '0' and StoredData = "010100001111" then SHout <= '1' after delay1 + 1295*delay_incr;
elsif nramp = '0' and StoredData = "010100010000" then SHout <= '1' after delay1 + 1296*delay_incr;
elsif nramp = '0' and StoredData = "010100010001" then SHout <= '1' after delay1 + 1297*delay_incr;
elsif nramp = '0' and StoredData = "010100010010" then SHout <= '1' after delay1 + 1298*delay_incr;
elsif nramp = '0' and StoredData = "010100010011" then SHout <= '1' after delay1 + 1299*delay_incr;
elsif nramp = '0' and StoredData = "010100010100" then SHout <= '1' after delay1 + 1300*delay_incr;
elsif nramp = '0' and StoredData = "010100010101" then SHout <= '1' after delay1 + 1301*delay_incr;
elsif nramp = '0' and StoredData = "010100010110" then SHout <= '1' after delay1 + 1302*delay_incr;
elsif nramp = '0' and StoredData = "010100010111" then SHout <= '1' after delay1 + 1303*delay_incr;
elsif nramp = '0' and StoredData = "010100011000" then SHout <= '1' after delay1 + 1304*delay_incr;
elsif nramp = '0' and StoredData = "010100011001" then SHout <= '1' after delay1 + 1305*delay_incr;
elsif nramp = '0' and StoredData = "010100011010" then SHout <= '1' after delay1 + 1306*delay_incr;
elsif nramp = '0' and StoredData = "010100011011" then SHout <= '1' after delay1 + 1307*delay_incr;
elsif nramp = '0' and StoredData = "010100011100" then SHout <= '1' after delay1 + 1308*delay_incr;
elsif nramp = '0' and StoredData = "010100011101" then SHout <= '1' after delay1 + 1309*delay_incr;
elsif nramp = '0' and StoredData = "010100011110" then SHout <= '1' after delay1 + 1310*delay_incr;
elsif nramp = '0' and StoredData = "010100011111" then SHout <= '1' after delay1 + 1311*delay_incr;
elsif nramp = '0' and StoredData = "010100100000" then SHout <= '1' after delay1 + 1312*delay_incr;
elsif nramp = '0' and StoredData = "010100100001" then SHout <= '1' after delay1 + 1313*delay_incr;
elsif nramp = '0' and StoredData = "010100100010" then SHout <= '1' after delay1 + 1314*delay_incr;
elsif nramp = '0' and StoredData = "010100100011" then SHout <= '1' after delay1 + 1315*delay_incr;
elsif nramp = '0' and StoredData = "010100100100" then SHout <= '1' after delay1 + 1316*delay_incr;
elsif nramp = '0' and StoredData = "010100100101" then SHout <= '1' after delay1 + 1317*delay_incr;
elsif nramp = '0' and StoredData = "010100100110" then SHout <= '1' after delay1 + 1318*delay_incr;
elsif nramp = '0' and StoredData = "010100100111" then SHout <= '1' after delay1 + 1319*delay_incr;
elsif nramp = '0' and StoredData = "010100101000" then SHout <= '1' after delay1 + 1320*delay_incr;
elsif nramp = '0' and StoredData = "010100101001" then SHout <= '1' after delay1 + 1321*delay_incr;
elsif nramp = '0' and StoredData = "010100101010" then SHout <= '1' after delay1 + 1322*delay_incr;
elsif nramp = '0' and StoredData = "010100101011" then SHout <= '1' after delay1 + 1323*delay_incr;
elsif nramp = '0' and StoredData = "010100101100" then SHout <= '1' after delay1 + 1324*delay_incr;
elsif nramp = '0' and StoredData = "010100101101" then SHout <= '1' after delay1 + 1325*delay_incr;
elsif nramp = '0' and StoredData = "010100101110" then SHout <= '1' after delay1 + 1326*delay_incr;
elsif nramp = '0' and StoredData = "010100101111" then SHout <= '1' after delay1 + 1327*delay_incr;
elsif nramp = '0' and StoredData = "010100110000" then SHout <= '1' after delay1 + 1328*delay_incr;
elsif nramp = '0' and StoredData = "010100110001" then SHout <= '1' after delay1 + 1329*delay_incr;
elsif nramp = '0' and StoredData = "010100110010" then SHout <= '1' after delay1 + 1330*delay_incr;
elsif nramp = '0' and StoredData = "010100110011" then SHout <= '1' after delay1 + 1331*delay_incr;
elsif nramp = '0' and StoredData = "010100110100" then SHout <= '1' after delay1 + 1332*delay_incr;
elsif nramp = '0' and StoredData = "010100110101" then SHout <= '1' after delay1 + 1333*delay_incr;
elsif nramp = '0' and StoredData = "010100110110" then SHout <= '1' after delay1 + 1334*delay_incr;
elsif nramp = '0' and StoredData = "010100110111" then SHout <= '1' after delay1 + 1335*delay_incr;
elsif nramp = '0' and StoredData = "010100111000" then SHout <= '1' after delay1 + 1336*delay_incr;
elsif nramp = '0' and StoredData = "010100111001" then SHout <= '1' after delay1 + 1337*delay_incr;
elsif nramp = '0' and StoredData = "010100111010" then SHout <= '1' after delay1 + 1338*delay_incr;
elsif nramp = '0' and StoredData = "010100111011" then SHout <= '1' after delay1 + 1339*delay_incr;
elsif nramp = '0' and StoredData = "010100111100" then SHout <= '1' after delay1 + 1340*delay_incr;
elsif nramp = '0' and StoredData = "010100111101" then SHout <= '1' after delay1 + 1341*delay_incr;
elsif nramp = '0' and StoredData = "010100111110" then SHout <= '1' after delay1 + 1342*delay_incr;
elsif nramp = '0' and StoredData = "010100111111" then SHout <= '1' after delay1 + 1343*delay_incr;
elsif nramp = '0' and StoredData = "010101000000" then SHout <= '1' after delay1 + 1344*delay_incr;
elsif nramp = '0' and StoredData = "010101000001" then SHout <= '1' after delay1 + 1345*delay_incr;
elsif nramp = '0' and StoredData = "010101000010" then SHout <= '1' after delay1 + 1346*delay_incr;
elsif nramp = '0' and StoredData = "010101000011" then SHout <= '1' after delay1 + 1347*delay_incr;
elsif nramp = '0' and StoredData = "010101000100" then SHout <= '1' after delay1 + 1348*delay_incr;
elsif nramp = '0' and StoredData = "010101000101" then SHout <= '1' after delay1 + 1349*delay_incr;
elsif nramp = '0' and StoredData = "010101000110" then SHout <= '1' after delay1 + 1350*delay_incr;
elsif nramp = '0' and StoredData = "010101000111" then SHout <= '1' after delay1 + 1351*delay_incr;
elsif nramp = '0' and StoredData = "010101001000" then SHout <= '1' after delay1 + 1352*delay_incr;
elsif nramp = '0' and StoredData = "010101001001" then SHout <= '1' after delay1 + 1353*delay_incr;
elsif nramp = '0' and StoredData = "010101001010" then SHout <= '1' after delay1 + 1354*delay_incr;
elsif nramp = '0' and StoredData = "010101001011" then SHout <= '1' after delay1 + 1355*delay_incr;
elsif nramp = '0' and StoredData = "010101001100" then SHout <= '1' after delay1 + 1356*delay_incr;
elsif nramp = '0' and StoredData = "010101001101" then SHout <= '1' after delay1 + 1357*delay_incr;
elsif nramp = '0' and StoredData = "010101001110" then SHout <= '1' after delay1 + 1358*delay_incr;
elsif nramp = '0' and StoredData = "010101001111" then SHout <= '1' after delay1 + 1359*delay_incr;
elsif nramp = '0' and StoredData = "010101010000" then SHout <= '1' after delay1 + 1360*delay_incr;
elsif nramp = '0' and StoredData = "010101010001" then SHout <= '1' after delay1 + 1361*delay_incr;
elsif nramp = '0' and StoredData = "010101010010" then SHout <= '1' after delay1 + 1362*delay_incr;
elsif nramp = '0' and StoredData = "010101010011" then SHout <= '1' after delay1 + 1363*delay_incr;
elsif nramp = '0' and StoredData = "010101010100" then SHout <= '1' after delay1 + 1364*delay_incr;
elsif nramp = '0' and StoredData = "010101010101" then SHout <= '1' after delay1 + 1365*delay_incr;
elsif nramp = '0' and StoredData = "010101010110" then SHout <= '1' after delay1 + 1366*delay_incr;
elsif nramp = '0' and StoredData = "010101010111" then SHout <= '1' after delay1 + 1367*delay_incr;
elsif nramp = '0' and StoredData = "010101011000" then SHout <= '1' after delay1 + 1368*delay_incr;
elsif nramp = '0' and StoredData = "010101011001" then SHout <= '1' after delay1 + 1369*delay_incr;
elsif nramp = '0' and StoredData = "010101011010" then SHout <= '1' after delay1 + 1370*delay_incr;
elsif nramp = '0' and StoredData = "010101011011" then SHout <= '1' after delay1 + 1371*delay_incr;
elsif nramp = '0' and StoredData = "010101011100" then SHout <= '1' after delay1 + 1372*delay_incr;
elsif nramp = '0' and StoredData = "010101011101" then SHout <= '1' after delay1 + 1373*delay_incr;
elsif nramp = '0' and StoredData = "010101011110" then SHout <= '1' after delay1 + 1374*delay_incr;
elsif nramp = '0' and StoredData = "010101011111" then SHout <= '1' after delay1 + 1375*delay_incr;
elsif nramp = '0' and StoredData = "010101100000" then SHout <= '1' after delay1 + 1376*delay_incr;
elsif nramp = '0' and StoredData = "010101100001" then SHout <= '1' after delay1 + 1377*delay_incr;
elsif nramp = '0' and StoredData = "010101100010" then SHout <= '1' after delay1 + 1378*delay_incr;
elsif nramp = '0' and StoredData = "010101100011" then SHout <= '1' after delay1 + 1379*delay_incr;
elsif nramp = '0' and StoredData = "010101100100" then SHout <= '1' after delay1 + 1380*delay_incr;
elsif nramp = '0' and StoredData = "010101100101" then SHout <= '1' after delay1 + 1381*delay_incr;
elsif nramp = '0' and StoredData = "010101100110" then SHout <= '1' after delay1 + 1382*delay_incr;
elsif nramp = '0' and StoredData = "010101100111" then SHout <= '1' after delay1 + 1383*delay_incr;
elsif nramp = '0' and StoredData = "010101101000" then SHout <= '1' after delay1 + 1384*delay_incr;
elsif nramp = '0' and StoredData = "010101101001" then SHout <= '1' after delay1 + 1385*delay_incr;
elsif nramp = '0' and StoredData = "010101101010" then SHout <= '1' after delay1 + 1386*delay_incr;
elsif nramp = '0' and StoredData = "010101101011" then SHout <= '1' after delay1 + 1387*delay_incr;
elsif nramp = '0' and StoredData = "010101101100" then SHout <= '1' after delay1 + 1388*delay_incr;
elsif nramp = '0' and StoredData = "010101101101" then SHout <= '1' after delay1 + 1389*delay_incr;
elsif nramp = '0' and StoredData = "010101101110" then SHout <= '1' after delay1 + 1390*delay_incr;
elsif nramp = '0' and StoredData = "010101101111" then SHout <= '1' after delay1 + 1391*delay_incr;
elsif nramp = '0' and StoredData = "010101110000" then SHout <= '1' after delay1 + 1392*delay_incr;
elsif nramp = '0' and StoredData = "010101110001" then SHout <= '1' after delay1 + 1393*delay_incr;
elsif nramp = '0' and StoredData = "010101110010" then SHout <= '1' after delay1 + 1394*delay_incr;
elsif nramp = '0' and StoredData = "010101110011" then SHout <= '1' after delay1 + 1395*delay_incr;
elsif nramp = '0' and StoredData = "010101110100" then SHout <= '1' after delay1 + 1396*delay_incr;
elsif nramp = '0' and StoredData = "010101110101" then SHout <= '1' after delay1 + 1397*delay_incr;
elsif nramp = '0' and StoredData = "010101110110" then SHout <= '1' after delay1 + 1398*delay_incr;
elsif nramp = '0' and StoredData = "010101110111" then SHout <= '1' after delay1 + 1399*delay_incr;
elsif nramp = '0' and StoredData = "010101111000" then SHout <= '1' after delay1 + 1400*delay_incr;
elsif nramp = '0' and StoredData = "010101111001" then SHout <= '1' after delay1 + 1401*delay_incr;
elsif nramp = '0' and StoredData = "010101111010" then SHout <= '1' after delay1 + 1402*delay_incr;
elsif nramp = '0' and StoredData = "010101111011" then SHout <= '1' after delay1 + 1403*delay_incr;
elsif nramp = '0' and StoredData = "010101111100" then SHout <= '1' after delay1 + 1404*delay_incr;
elsif nramp = '0' and StoredData = "010101111101" then SHout <= '1' after delay1 + 1405*delay_incr;
elsif nramp = '0' and StoredData = "010101111110" then SHout <= '1' after delay1 + 1406*delay_incr;
elsif nramp = '0' and StoredData = "010101111111" then SHout <= '1' after delay1 + 1407*delay_incr;
elsif nramp = '0' and StoredData = "010110000000" then SHout <= '1' after delay1 + 1408*delay_incr;
elsif nramp = '0' and StoredData = "010110000001" then SHout <= '1' after delay1 + 1409*delay_incr;
elsif nramp = '0' and StoredData = "010110000010" then SHout <= '1' after delay1 + 1410*delay_incr;
elsif nramp = '0' and StoredData = "010110000011" then SHout <= '1' after delay1 + 1411*delay_incr;
elsif nramp = '0' and StoredData = "010110000100" then SHout <= '1' after delay1 + 1412*delay_incr;
elsif nramp = '0' and StoredData = "010110000101" then SHout <= '1' after delay1 + 1413*delay_incr;
elsif nramp = '0' and StoredData = "010110000110" then SHout <= '1' after delay1 + 1414*delay_incr;
elsif nramp = '0' and StoredData = "010110000111" then SHout <= '1' after delay1 + 1415*delay_incr;
elsif nramp = '0' and StoredData = "010110001000" then SHout <= '1' after delay1 + 1416*delay_incr;
elsif nramp = '0' and StoredData = "010110001001" then SHout <= '1' after delay1 + 1417*delay_incr;
elsif nramp = '0' and StoredData = "010110001010" then SHout <= '1' after delay1 + 1418*delay_incr;
elsif nramp = '0' and StoredData = "010110001011" then SHout <= '1' after delay1 + 1419*delay_incr;
elsif nramp = '0' and StoredData = "010110001100" then SHout <= '1' after delay1 + 1420*delay_incr;
elsif nramp = '0' and StoredData = "010110001101" then SHout <= '1' after delay1 + 1421*delay_incr;
elsif nramp = '0' and StoredData = "010110001110" then SHout <= '1' after delay1 + 1422*delay_incr;
elsif nramp = '0' and StoredData = "010110001111" then SHout <= '1' after delay1 + 1423*delay_incr;
elsif nramp = '0' and StoredData = "010110010000" then SHout <= '1' after delay1 + 1424*delay_incr;
elsif nramp = '0' and StoredData = "010110010001" then SHout <= '1' after delay1 + 1425*delay_incr;
elsif nramp = '0' and StoredData = "010110010010" then SHout <= '1' after delay1 + 1426*delay_incr;
elsif nramp = '0' and StoredData = "010110010011" then SHout <= '1' after delay1 + 1427*delay_incr;
elsif nramp = '0' and StoredData = "010110010100" then SHout <= '1' after delay1 + 1428*delay_incr;
elsif nramp = '0' and StoredData = "010110010101" then SHout <= '1' after delay1 + 1429*delay_incr;
elsif nramp = '0' and StoredData = "010110010110" then SHout <= '1' after delay1 + 1430*delay_incr;
elsif nramp = '0' and StoredData = "010110010111" then SHout <= '1' after delay1 + 1431*delay_incr;
elsif nramp = '0' and StoredData = "010110011000" then SHout <= '1' after delay1 + 1432*delay_incr;
elsif nramp = '0' and StoredData = "010110011001" then SHout <= '1' after delay1 + 1433*delay_incr;
elsif nramp = '0' and StoredData = "010110011010" then SHout <= '1' after delay1 + 1434*delay_incr;
elsif nramp = '0' and StoredData = "010110011011" then SHout <= '1' after delay1 + 1435*delay_incr;
elsif nramp = '0' and StoredData = "010110011100" then SHout <= '1' after delay1 + 1436*delay_incr;
elsif nramp = '0' and StoredData = "010110011101" then SHout <= '1' after delay1 + 1437*delay_incr;
elsif nramp = '0' and StoredData = "010110011110" then SHout <= '1' after delay1 + 1438*delay_incr;
elsif nramp = '0' and StoredData = "010110011111" then SHout <= '1' after delay1 + 1439*delay_incr;
elsif nramp = '0' and StoredData = "010110100000" then SHout <= '1' after delay1 + 1440*delay_incr;
elsif nramp = '0' and StoredData = "010110100001" then SHout <= '1' after delay1 + 1441*delay_incr;
elsif nramp = '0' and StoredData = "010110100010" then SHout <= '1' after delay1 + 1442*delay_incr;
elsif nramp = '0' and StoredData = "010110100011" then SHout <= '1' after delay1 + 1443*delay_incr;
elsif nramp = '0' and StoredData = "010110100100" then SHout <= '1' after delay1 + 1444*delay_incr;
elsif nramp = '0' and StoredData = "010110100101" then SHout <= '1' after delay1 + 1445*delay_incr;
elsif nramp = '0' and StoredData = "010110100110" then SHout <= '1' after delay1 + 1446*delay_incr;
elsif nramp = '0' and StoredData = "010110100111" then SHout <= '1' after delay1 + 1447*delay_incr;
elsif nramp = '0' and StoredData = "010110101000" then SHout <= '1' after delay1 + 1448*delay_incr;
elsif nramp = '0' and StoredData = "010110101001" then SHout <= '1' after delay1 + 1449*delay_incr;
elsif nramp = '0' and StoredData = "010110101010" then SHout <= '1' after delay1 + 1450*delay_incr;
elsif nramp = '0' and StoredData = "010110101011" then SHout <= '1' after delay1 + 1451*delay_incr;
elsif nramp = '0' and StoredData = "010110101100" then SHout <= '1' after delay1 + 1452*delay_incr;
elsif nramp = '0' and StoredData = "010110101101" then SHout <= '1' after delay1 + 1453*delay_incr;
elsif nramp = '0' and StoredData = "010110101110" then SHout <= '1' after delay1 + 1454*delay_incr;
elsif nramp = '0' and StoredData = "010110101111" then SHout <= '1' after delay1 + 1455*delay_incr;
elsif nramp = '0' and StoredData = "010110110000" then SHout <= '1' after delay1 + 1456*delay_incr;
elsif nramp = '0' and StoredData = "010110110001" then SHout <= '1' after delay1 + 1457*delay_incr;
elsif nramp = '0' and StoredData = "010110110010" then SHout <= '1' after delay1 + 1458*delay_incr;
elsif nramp = '0' and StoredData = "010110110011" then SHout <= '1' after delay1 + 1459*delay_incr;
elsif nramp = '0' and StoredData = "010110110100" then SHout <= '1' after delay1 + 1460*delay_incr;
elsif nramp = '0' and StoredData = "010110110101" then SHout <= '1' after delay1 + 1461*delay_incr;
elsif nramp = '0' and StoredData = "010110110110" then SHout <= '1' after delay1 + 1462*delay_incr;
elsif nramp = '0' and StoredData = "010110110111" then SHout <= '1' after delay1 + 1463*delay_incr;
elsif nramp = '0' and StoredData = "010110111000" then SHout <= '1' after delay1 + 1464*delay_incr;
elsif nramp = '0' and StoredData = "010110111001" then SHout <= '1' after delay1 + 1465*delay_incr;
elsif nramp = '0' and StoredData = "010110111010" then SHout <= '1' after delay1 + 1466*delay_incr;
elsif nramp = '0' and StoredData = "010110111011" then SHout <= '1' after delay1 + 1467*delay_incr;
elsif nramp = '0' and StoredData = "010110111100" then SHout <= '1' after delay1 + 1468*delay_incr;
elsif nramp = '0' and StoredData = "010110111101" then SHout <= '1' after delay1 + 1469*delay_incr;
elsif nramp = '0' and StoredData = "010110111110" then SHout <= '1' after delay1 + 1470*delay_incr;
elsif nramp = '0' and StoredData = "010110111111" then SHout <= '1' after delay1 + 1471*delay_incr;
elsif nramp = '0' and StoredData = "010111000000" then SHout <= '1' after delay1 + 1472*delay_incr;
elsif nramp = '0' and StoredData = "010111000001" then SHout <= '1' after delay1 + 1473*delay_incr;
elsif nramp = '0' and StoredData = "010111000010" then SHout <= '1' after delay1 + 1474*delay_incr;
elsif nramp = '0' and StoredData = "010111000011" then SHout <= '1' after delay1 + 1475*delay_incr;
elsif nramp = '0' and StoredData = "010111000100" then SHout <= '1' after delay1 + 1476*delay_incr;
elsif nramp = '0' and StoredData = "010111000101" then SHout <= '1' after delay1 + 1477*delay_incr;
elsif nramp = '0' and StoredData = "010111000110" then SHout <= '1' after delay1 + 1478*delay_incr;
elsif nramp = '0' and StoredData = "010111000111" then SHout <= '1' after delay1 + 1479*delay_incr;
elsif nramp = '0' and StoredData = "010111001000" then SHout <= '1' after delay1 + 1480*delay_incr;
elsif nramp = '0' and StoredData = "010111001001" then SHout <= '1' after delay1 + 1481*delay_incr;
elsif nramp = '0' and StoredData = "010111001010" then SHout <= '1' after delay1 + 1482*delay_incr;
elsif nramp = '0' and StoredData = "010111001011" then SHout <= '1' after delay1 + 1483*delay_incr;
elsif nramp = '0' and StoredData = "010111001100" then SHout <= '1' after delay1 + 1484*delay_incr;
elsif nramp = '0' and StoredData = "010111001101" then SHout <= '1' after delay1 + 1485*delay_incr;
elsif nramp = '0' and StoredData = "010111001110" then SHout <= '1' after delay1 + 1486*delay_incr;
elsif nramp = '0' and StoredData = "010111001111" then SHout <= '1' after delay1 + 1487*delay_incr;
elsif nramp = '0' and StoredData = "010111010000" then SHout <= '1' after delay1 + 1488*delay_incr;
elsif nramp = '0' and StoredData = "010111010001" then SHout <= '1' after delay1 + 1489*delay_incr;
elsif nramp = '0' and StoredData = "010111010010" then SHout <= '1' after delay1 + 1490*delay_incr;
elsif nramp = '0' and StoredData = "010111010011" then SHout <= '1' after delay1 + 1491*delay_incr;
elsif nramp = '0' and StoredData = "010111010100" then SHout <= '1' after delay1 + 1492*delay_incr;
elsif nramp = '0' and StoredData = "010111010101" then SHout <= '1' after delay1 + 1493*delay_incr;
elsif nramp = '0' and StoredData = "010111010110" then SHout <= '1' after delay1 + 1494*delay_incr;
elsif nramp = '0' and StoredData = "010111010111" then SHout <= '1' after delay1 + 1495*delay_incr;
elsif nramp = '0' and StoredData = "010111011000" then SHout <= '1' after delay1 + 1496*delay_incr;
elsif nramp = '0' and StoredData = "010111011001" then SHout <= '1' after delay1 + 1497*delay_incr;
elsif nramp = '0' and StoredData = "010111011010" then SHout <= '1' after delay1 + 1498*delay_incr;
elsif nramp = '0' and StoredData = "010111011011" then SHout <= '1' after delay1 + 1499*delay_incr;
elsif nramp = '0' and StoredData = "010111011100" then SHout <= '1' after delay1 + 1500*delay_incr;
elsif nramp = '0' and StoredData = "010111011101" then SHout <= '1' after delay1 + 1501*delay_incr;
elsif nramp = '0' and StoredData = "010111011110" then SHout <= '1' after delay1 + 1502*delay_incr;
elsif nramp = '0' and StoredData = "010111011111" then SHout <= '1' after delay1 + 1503*delay_incr;
elsif nramp = '0' and StoredData = "010111100000" then SHout <= '1' after delay1 + 1504*delay_incr;
elsif nramp = '0' and StoredData = "010111100001" then SHout <= '1' after delay1 + 1505*delay_incr;
elsif nramp = '0' and StoredData = "010111100010" then SHout <= '1' after delay1 + 1506*delay_incr;
elsif nramp = '0' and StoredData = "010111100011" then SHout <= '1' after delay1 + 1507*delay_incr;
elsif nramp = '0' and StoredData = "010111100100" then SHout <= '1' after delay1 + 1508*delay_incr;
elsif nramp = '0' and StoredData = "010111100101" then SHout <= '1' after delay1 + 1509*delay_incr;
elsif nramp = '0' and StoredData = "010111100110" then SHout <= '1' after delay1 + 1510*delay_incr;
elsif nramp = '0' and StoredData = "010111100111" then SHout <= '1' after delay1 + 1511*delay_incr;
elsif nramp = '0' and StoredData = "010111101000" then SHout <= '1' after delay1 + 1512*delay_incr;
elsif nramp = '0' and StoredData = "010111101001" then SHout <= '1' after delay1 + 1513*delay_incr;
elsif nramp = '0' and StoredData = "010111101010" then SHout <= '1' after delay1 + 1514*delay_incr;
elsif nramp = '0' and StoredData = "010111101011" then SHout <= '1' after delay1 + 1515*delay_incr;
elsif nramp = '0' and StoredData = "010111101100" then SHout <= '1' after delay1 + 1516*delay_incr;
elsif nramp = '0' and StoredData = "010111101101" then SHout <= '1' after delay1 + 1517*delay_incr;
elsif nramp = '0' and StoredData = "010111101110" then SHout <= '1' after delay1 + 1518*delay_incr;
elsif nramp = '0' and StoredData = "010111101111" then SHout <= '1' after delay1 + 1519*delay_incr;
elsif nramp = '0' and StoredData = "010111110000" then SHout <= '1' after delay1 + 1520*delay_incr;
elsif nramp = '0' and StoredData = "010111110001" then SHout <= '1' after delay1 + 1521*delay_incr;
elsif nramp = '0' and StoredData = "010111110010" then SHout <= '1' after delay1 + 1522*delay_incr;
elsif nramp = '0' and StoredData = "010111110011" then SHout <= '1' after delay1 + 1523*delay_incr;
elsif nramp = '0' and StoredData = "010111110100" then SHout <= '1' after delay1 + 1524*delay_incr;
elsif nramp = '0' and StoredData = "010111110101" then SHout <= '1' after delay1 + 1525*delay_incr;
elsif nramp = '0' and StoredData = "010111110110" then SHout <= '1' after delay1 + 1526*delay_incr;
elsif nramp = '0' and StoredData = "010111110111" then SHout <= '1' after delay1 + 1527*delay_incr;
elsif nramp = '0' and StoredData = "010111111000" then SHout <= '1' after delay1 + 1528*delay_incr;
elsif nramp = '0' and StoredData = "010111111001" then SHout <= '1' after delay1 + 1529*delay_incr;
elsif nramp = '0' and StoredData = "010111111010" then SHout <= '1' after delay1 + 1530*delay_incr;
elsif nramp = '0' and StoredData = "010111111011" then SHout <= '1' after delay1 + 1531*delay_incr;
elsif nramp = '0' and StoredData = "010111111100" then SHout <= '1' after delay1 + 1532*delay_incr;
elsif nramp = '0' and StoredData = "010111111101" then SHout <= '1' after delay1 + 1533*delay_incr;
elsif nramp = '0' and StoredData = "010111111110" then SHout <= '1' after delay1 + 1534*delay_incr;
elsif nramp = '0' and StoredData = "010111111111" then SHout <= '1' after delay1 + 1535*delay_incr;
elsif nramp = '0' and StoredData = "011000000000" then SHout <= '1' after delay1 + 1536*delay_incr;
elsif nramp = '0' and StoredData = "011000000001" then SHout <= '1' after delay1 + 1537*delay_incr;
elsif nramp = '0' and StoredData = "011000000010" then SHout <= '1' after delay1 + 1538*delay_incr;
elsif nramp = '0' and StoredData = "011000000011" then SHout <= '1' after delay1 + 1539*delay_incr;
elsif nramp = '0' and StoredData = "011000000100" then SHout <= '1' after delay1 + 1540*delay_incr;
elsif nramp = '0' and StoredData = "011000000101" then SHout <= '1' after delay1 + 1541*delay_incr;
elsif nramp = '0' and StoredData = "011000000110" then SHout <= '1' after delay1 + 1542*delay_incr;
elsif nramp = '0' and StoredData = "011000000111" then SHout <= '1' after delay1 + 1543*delay_incr;
elsif nramp = '0' and StoredData = "011000001000" then SHout <= '1' after delay1 + 1544*delay_incr;
elsif nramp = '0' and StoredData = "011000001001" then SHout <= '1' after delay1 + 1545*delay_incr;
elsif nramp = '0' and StoredData = "011000001010" then SHout <= '1' after delay1 + 1546*delay_incr;
elsif nramp = '0' and StoredData = "011000001011" then SHout <= '1' after delay1 + 1547*delay_incr;
elsif nramp = '0' and StoredData = "011000001100" then SHout <= '1' after delay1 + 1548*delay_incr;
elsif nramp = '0' and StoredData = "011000001101" then SHout <= '1' after delay1 + 1549*delay_incr;
elsif nramp = '0' and StoredData = "011000001110" then SHout <= '1' after delay1 + 1550*delay_incr;
elsif nramp = '0' and StoredData = "011000001111" then SHout <= '1' after delay1 + 1551*delay_incr;
elsif nramp = '0' and StoredData = "011000010000" then SHout <= '1' after delay1 + 1552*delay_incr;
elsif nramp = '0' and StoredData = "011000010001" then SHout <= '1' after delay1 + 1553*delay_incr;
elsif nramp = '0' and StoredData = "011000010010" then SHout <= '1' after delay1 + 1554*delay_incr;
elsif nramp = '0' and StoredData = "011000010011" then SHout <= '1' after delay1 + 1555*delay_incr;
elsif nramp = '0' and StoredData = "011000010100" then SHout <= '1' after delay1 + 1556*delay_incr;
elsif nramp = '0' and StoredData = "011000010101" then SHout <= '1' after delay1 + 1557*delay_incr;
elsif nramp = '0' and StoredData = "011000010110" then SHout <= '1' after delay1 + 1558*delay_incr;
elsif nramp = '0' and StoredData = "011000010111" then SHout <= '1' after delay1 + 1559*delay_incr;
elsif nramp = '0' and StoredData = "011000011000" then SHout <= '1' after delay1 + 1560*delay_incr;
elsif nramp = '0' and StoredData = "011000011001" then SHout <= '1' after delay1 + 1561*delay_incr;
elsif nramp = '0' and StoredData = "011000011010" then SHout <= '1' after delay1 + 1562*delay_incr;
elsif nramp = '0' and StoredData = "011000011011" then SHout <= '1' after delay1 + 1563*delay_incr;
elsif nramp = '0' and StoredData = "011000011100" then SHout <= '1' after delay1 + 1564*delay_incr;
elsif nramp = '0' and StoredData = "011000011101" then SHout <= '1' after delay1 + 1565*delay_incr;
elsif nramp = '0' and StoredData = "011000011110" then SHout <= '1' after delay1 + 1566*delay_incr;
elsif nramp = '0' and StoredData = "011000011111" then SHout <= '1' after delay1 + 1567*delay_incr;
elsif nramp = '0' and StoredData = "011000100000" then SHout <= '1' after delay1 + 1568*delay_incr;
elsif nramp = '0' and StoredData = "011000100001" then SHout <= '1' after delay1 + 1569*delay_incr;
elsif nramp = '0' and StoredData = "011000100010" then SHout <= '1' after delay1 + 1570*delay_incr;
elsif nramp = '0' and StoredData = "011000100011" then SHout <= '1' after delay1 + 1571*delay_incr;
elsif nramp = '0' and StoredData = "011000100100" then SHout <= '1' after delay1 + 1572*delay_incr;
elsif nramp = '0' and StoredData = "011000100101" then SHout <= '1' after delay1 + 1573*delay_incr;
elsif nramp = '0' and StoredData = "011000100110" then SHout <= '1' after delay1 + 1574*delay_incr;
elsif nramp = '0' and StoredData = "011000100111" then SHout <= '1' after delay1 + 1575*delay_incr;
elsif nramp = '0' and StoredData = "011000101000" then SHout <= '1' after delay1 + 1576*delay_incr;
elsif nramp = '0' and StoredData = "011000101001" then SHout <= '1' after delay1 + 1577*delay_incr;
elsif nramp = '0' and StoredData = "011000101010" then SHout <= '1' after delay1 + 1578*delay_incr;
elsif nramp = '0' and StoredData = "011000101011" then SHout <= '1' after delay1 + 1579*delay_incr;
elsif nramp = '0' and StoredData = "011000101100" then SHout <= '1' after delay1 + 1580*delay_incr;
elsif nramp = '0' and StoredData = "011000101101" then SHout <= '1' after delay1 + 1581*delay_incr;
elsif nramp = '0' and StoredData = "011000101110" then SHout <= '1' after delay1 + 1582*delay_incr;
elsif nramp = '0' and StoredData = "011000101111" then SHout <= '1' after delay1 + 1583*delay_incr;
elsif nramp = '0' and StoredData = "011000110000" then SHout <= '1' after delay1 + 1584*delay_incr;
elsif nramp = '0' and StoredData = "011000110001" then SHout <= '1' after delay1 + 1585*delay_incr;
elsif nramp = '0' and StoredData = "011000110010" then SHout <= '1' after delay1 + 1586*delay_incr;
elsif nramp = '0' and StoredData = "011000110011" then SHout <= '1' after delay1 + 1587*delay_incr;
elsif nramp = '0' and StoredData = "011000110100" then SHout <= '1' after delay1 + 1588*delay_incr;
elsif nramp = '0' and StoredData = "011000110101" then SHout <= '1' after delay1 + 1589*delay_incr;
elsif nramp = '0' and StoredData = "011000110110" then SHout <= '1' after delay1 + 1590*delay_incr;
elsif nramp = '0' and StoredData = "011000110111" then SHout <= '1' after delay1 + 1591*delay_incr;
elsif nramp = '0' and StoredData = "011000111000" then SHout <= '1' after delay1 + 1592*delay_incr;
elsif nramp = '0' and StoredData = "011000111001" then SHout <= '1' after delay1 + 1593*delay_incr;
elsif nramp = '0' and StoredData = "011000111010" then SHout <= '1' after delay1 + 1594*delay_incr;
elsif nramp = '0' and StoredData = "011000111011" then SHout <= '1' after delay1 + 1595*delay_incr;
elsif nramp = '0' and StoredData = "011000111100" then SHout <= '1' after delay1 + 1596*delay_incr;
elsif nramp = '0' and StoredData = "011000111101" then SHout <= '1' after delay1 + 1597*delay_incr;
elsif nramp = '0' and StoredData = "011000111110" then SHout <= '1' after delay1 + 1598*delay_incr;
elsif nramp = '0' and StoredData = "011000111111" then SHout <= '1' after delay1 + 1599*delay_incr;
elsif nramp = '0' and StoredData = "011001000000" then SHout <= '1' after delay1 + 1600*delay_incr;
elsif nramp = '0' and StoredData = "011001000001" then SHout <= '1' after delay1 + 1601*delay_incr;
elsif nramp = '0' and StoredData = "011001000010" then SHout <= '1' after delay1 + 1602*delay_incr;
elsif nramp = '0' and StoredData = "011001000011" then SHout <= '1' after delay1 + 1603*delay_incr;
elsif nramp = '0' and StoredData = "011001000100" then SHout <= '1' after delay1 + 1604*delay_incr;
elsif nramp = '0' and StoredData = "011001000101" then SHout <= '1' after delay1 + 1605*delay_incr;
elsif nramp = '0' and StoredData = "011001000110" then SHout <= '1' after delay1 + 1606*delay_incr;
elsif nramp = '0' and StoredData = "011001000111" then SHout <= '1' after delay1 + 1607*delay_incr;
elsif nramp = '0' and StoredData = "011001001000" then SHout <= '1' after delay1 + 1608*delay_incr;
elsif nramp = '0' and StoredData = "011001001001" then SHout <= '1' after delay1 + 1609*delay_incr;
elsif nramp = '0' and StoredData = "011001001010" then SHout <= '1' after delay1 + 1610*delay_incr;
elsif nramp = '0' and StoredData = "011001001011" then SHout <= '1' after delay1 + 1611*delay_incr;
elsif nramp = '0' and StoredData = "011001001100" then SHout <= '1' after delay1 + 1612*delay_incr;
elsif nramp = '0' and StoredData = "011001001101" then SHout <= '1' after delay1 + 1613*delay_incr;
elsif nramp = '0' and StoredData = "011001001110" then SHout <= '1' after delay1 + 1614*delay_incr;
elsif nramp = '0' and StoredData = "011001001111" then SHout <= '1' after delay1 + 1615*delay_incr;
elsif nramp = '0' and StoredData = "011001010000" then SHout <= '1' after delay1 + 1616*delay_incr;
elsif nramp = '0' and StoredData = "011001010001" then SHout <= '1' after delay1 + 1617*delay_incr;
elsif nramp = '0' and StoredData = "011001010010" then SHout <= '1' after delay1 + 1618*delay_incr;
elsif nramp = '0' and StoredData = "011001010011" then SHout <= '1' after delay1 + 1619*delay_incr;
elsif nramp = '0' and StoredData = "011001010100" then SHout <= '1' after delay1 + 1620*delay_incr;
elsif nramp = '0' and StoredData = "011001010101" then SHout <= '1' after delay1 + 1621*delay_incr;
elsif nramp = '0' and StoredData = "011001010110" then SHout <= '1' after delay1 + 1622*delay_incr;
elsif nramp = '0' and StoredData = "011001010111" then SHout <= '1' after delay1 + 1623*delay_incr;
elsif nramp = '0' and StoredData = "011001011000" then SHout <= '1' after delay1 + 1624*delay_incr;
elsif nramp = '0' and StoredData = "011001011001" then SHout <= '1' after delay1 + 1625*delay_incr;
elsif nramp = '0' and StoredData = "011001011010" then SHout <= '1' after delay1 + 1626*delay_incr;
elsif nramp = '0' and StoredData = "011001011011" then SHout <= '1' after delay1 + 1627*delay_incr;
elsif nramp = '0' and StoredData = "011001011100" then SHout <= '1' after delay1 + 1628*delay_incr;
elsif nramp = '0' and StoredData = "011001011101" then SHout <= '1' after delay1 + 1629*delay_incr;
elsif nramp = '0' and StoredData = "011001011110" then SHout <= '1' after delay1 + 1630*delay_incr;
elsif nramp = '0' and StoredData = "011001011111" then SHout <= '1' after delay1 + 1631*delay_incr;
elsif nramp = '0' and StoredData = "011001100000" then SHout <= '1' after delay1 + 1632*delay_incr;
elsif nramp = '0' and StoredData = "011001100001" then SHout <= '1' after delay1 + 1633*delay_incr;
elsif nramp = '0' and StoredData = "011001100010" then SHout <= '1' after delay1 + 1634*delay_incr;
elsif nramp = '0' and StoredData = "011001100011" then SHout <= '1' after delay1 + 1635*delay_incr;
elsif nramp = '0' and StoredData = "011001100100" then SHout <= '1' after delay1 + 1636*delay_incr;
elsif nramp = '0' and StoredData = "011001100101" then SHout <= '1' after delay1 + 1637*delay_incr;
elsif nramp = '0' and StoredData = "011001100110" then SHout <= '1' after delay1 + 1638*delay_incr;
elsif nramp = '0' and StoredData = "011001100111" then SHout <= '1' after delay1 + 1639*delay_incr;
elsif nramp = '0' and StoredData = "011001101000" then SHout <= '1' after delay1 + 1640*delay_incr;
elsif nramp = '0' and StoredData = "011001101001" then SHout <= '1' after delay1 + 1641*delay_incr;
elsif nramp = '0' and StoredData = "011001101010" then SHout <= '1' after delay1 + 1642*delay_incr;
elsif nramp = '0' and StoredData = "011001101011" then SHout <= '1' after delay1 + 1643*delay_incr;
elsif nramp = '0' and StoredData = "011001101100" then SHout <= '1' after delay1 + 1644*delay_incr;
elsif nramp = '0' and StoredData = "011001101101" then SHout <= '1' after delay1 + 1645*delay_incr;
elsif nramp = '0' and StoredData = "011001101110" then SHout <= '1' after delay1 + 1646*delay_incr;
elsif nramp = '0' and StoredData = "011001101111" then SHout <= '1' after delay1 + 1647*delay_incr;
elsif nramp = '0' and StoredData = "011001110000" then SHout <= '1' after delay1 + 1648*delay_incr;
elsif nramp = '0' and StoredData = "011001110001" then SHout <= '1' after delay1 + 1649*delay_incr;
elsif nramp = '0' and StoredData = "011001110010" then SHout <= '1' after delay1 + 1650*delay_incr;
elsif nramp = '0' and StoredData = "011001110011" then SHout <= '1' after delay1 + 1651*delay_incr;
elsif nramp = '0' and StoredData = "011001110100" then SHout <= '1' after delay1 + 1652*delay_incr;
elsif nramp = '0' and StoredData = "011001110101" then SHout <= '1' after delay1 + 1653*delay_incr;
elsif nramp = '0' and StoredData = "011001110110" then SHout <= '1' after delay1 + 1654*delay_incr;
elsif nramp = '0' and StoredData = "011001110111" then SHout <= '1' after delay1 + 1655*delay_incr;
elsif nramp = '0' and StoredData = "011001111000" then SHout <= '1' after delay1 + 1656*delay_incr;
elsif nramp = '0' and StoredData = "011001111001" then SHout <= '1' after delay1 + 1657*delay_incr;
elsif nramp = '0' and StoredData = "011001111010" then SHout <= '1' after delay1 + 1658*delay_incr;
elsif nramp = '0' and StoredData = "011001111011" then SHout <= '1' after delay1 + 1659*delay_incr;
elsif nramp = '0' and StoredData = "011001111100" then SHout <= '1' after delay1 + 1660*delay_incr;
elsif nramp = '0' and StoredData = "011001111101" then SHout <= '1' after delay1 + 1661*delay_incr;
elsif nramp = '0' and StoredData = "011001111110" then SHout <= '1' after delay1 + 1662*delay_incr;
elsif nramp = '0' and StoredData = "011001111111" then SHout <= '1' after delay1 + 1663*delay_incr;
elsif nramp = '0' and StoredData = "011010000000" then SHout <= '1' after delay1 + 1664*delay_incr;
elsif nramp = '0' and StoredData = "011010000001" then SHout <= '1' after delay1 + 1665*delay_incr;
elsif nramp = '0' and StoredData = "011010000010" then SHout <= '1' after delay1 + 1666*delay_incr;
elsif nramp = '0' and StoredData = "011010000011" then SHout <= '1' after delay1 + 1667*delay_incr;
elsif nramp = '0' and StoredData = "011010000100" then SHout <= '1' after delay1 + 1668*delay_incr;
elsif nramp = '0' and StoredData = "011010000101" then SHout <= '1' after delay1 + 1669*delay_incr;
elsif nramp = '0' and StoredData = "011010000110" then SHout <= '1' after delay1 + 1670*delay_incr;
elsif nramp = '0' and StoredData = "011010000111" then SHout <= '1' after delay1 + 1671*delay_incr;
elsif nramp = '0' and StoredData = "011010001000" then SHout <= '1' after delay1 + 1672*delay_incr;
elsif nramp = '0' and StoredData = "011010001001" then SHout <= '1' after delay1 + 1673*delay_incr;
elsif nramp = '0' and StoredData = "011010001010" then SHout <= '1' after delay1 + 1674*delay_incr;
elsif nramp = '0' and StoredData = "011010001011" then SHout <= '1' after delay1 + 1675*delay_incr;
elsif nramp = '0' and StoredData = "011010001100" then SHout <= '1' after delay1 + 1676*delay_incr;
elsif nramp = '0' and StoredData = "011010001101" then SHout <= '1' after delay1 + 1677*delay_incr;
elsif nramp = '0' and StoredData = "011010001110" then SHout <= '1' after delay1 + 1678*delay_incr;
elsif nramp = '0' and StoredData = "011010001111" then SHout <= '1' after delay1 + 1679*delay_incr;
elsif nramp = '0' and StoredData = "011010010000" then SHout <= '1' after delay1 + 1680*delay_incr;
elsif nramp = '0' and StoredData = "011010010001" then SHout <= '1' after delay1 + 1681*delay_incr;
elsif nramp = '0' and StoredData = "011010010010" then SHout <= '1' after delay1 + 1682*delay_incr;
elsif nramp = '0' and StoredData = "011010010011" then SHout <= '1' after delay1 + 1683*delay_incr;
elsif nramp = '0' and StoredData = "011010010100" then SHout <= '1' after delay1 + 1684*delay_incr;
elsif nramp = '0' and StoredData = "011010010101" then SHout <= '1' after delay1 + 1685*delay_incr;
elsif nramp = '0' and StoredData = "011010010110" then SHout <= '1' after delay1 + 1686*delay_incr;
elsif nramp = '0' and StoredData = "011010010111" then SHout <= '1' after delay1 + 1687*delay_incr;
elsif nramp = '0' and StoredData = "011010011000" then SHout <= '1' after delay1 + 1688*delay_incr;
elsif nramp = '0' and StoredData = "011010011001" then SHout <= '1' after delay1 + 1689*delay_incr;
elsif nramp = '0' and StoredData = "011010011010" then SHout <= '1' after delay1 + 1690*delay_incr;
elsif nramp = '0' and StoredData = "011010011011" then SHout <= '1' after delay1 + 1691*delay_incr;
elsif nramp = '0' and StoredData = "011010011100" then SHout <= '1' after delay1 + 1692*delay_incr;
elsif nramp = '0' and StoredData = "011010011101" then SHout <= '1' after delay1 + 1693*delay_incr;
elsif nramp = '0' and StoredData = "011010011110" then SHout <= '1' after delay1 + 1694*delay_incr;
elsif nramp = '0' and StoredData = "011010011111" then SHout <= '1' after delay1 + 1695*delay_incr;
elsif nramp = '0' and StoredData = "011010100000" then SHout <= '1' after delay1 + 1696*delay_incr;
elsif nramp = '0' and StoredData = "011010100001" then SHout <= '1' after delay1 + 1697*delay_incr;
elsif nramp = '0' and StoredData = "011010100010" then SHout <= '1' after delay1 + 1698*delay_incr;
elsif nramp = '0' and StoredData = "011010100011" then SHout <= '1' after delay1 + 1699*delay_incr;
elsif nramp = '0' and StoredData = "011010100100" then SHout <= '1' after delay1 + 1700*delay_incr;
elsif nramp = '0' and StoredData = "011010100101" then SHout <= '1' after delay1 + 1701*delay_incr;
elsif nramp = '0' and StoredData = "011010100110" then SHout <= '1' after delay1 + 1702*delay_incr;
elsif nramp = '0' and StoredData = "011010100111" then SHout <= '1' after delay1 + 1703*delay_incr;
elsif nramp = '0' and StoredData = "011010101000" then SHout <= '1' after delay1 + 1704*delay_incr;
elsif nramp = '0' and StoredData = "011010101001" then SHout <= '1' after delay1 + 1705*delay_incr;
elsif nramp = '0' and StoredData = "011010101010" then SHout <= '1' after delay1 + 1706*delay_incr;
elsif nramp = '0' and StoredData = "011010101011" then SHout <= '1' after delay1 + 1707*delay_incr;
elsif nramp = '0' and StoredData = "011010101100" then SHout <= '1' after delay1 + 1708*delay_incr;
elsif nramp = '0' and StoredData = "011010101101" then SHout <= '1' after delay1 + 1709*delay_incr;
elsif nramp = '0' and StoredData = "011010101110" then SHout <= '1' after delay1 + 1710*delay_incr;
elsif nramp = '0' and StoredData = "011010101111" then SHout <= '1' after delay1 + 1711*delay_incr;
elsif nramp = '0' and StoredData = "011010110000" then SHout <= '1' after delay1 + 1712*delay_incr;
elsif nramp = '0' and StoredData = "011010110001" then SHout <= '1' after delay1 + 1713*delay_incr;
elsif nramp = '0' and StoredData = "011010110010" then SHout <= '1' after delay1 + 1714*delay_incr;
elsif nramp = '0' and StoredData = "011010110011" then SHout <= '1' after delay1 + 1715*delay_incr;
elsif nramp = '0' and StoredData = "011010110100" then SHout <= '1' after delay1 + 1716*delay_incr;
elsif nramp = '0' and StoredData = "011010110101" then SHout <= '1' after delay1 + 1717*delay_incr;
elsif nramp = '0' and StoredData = "011010110110" then SHout <= '1' after delay1 + 1718*delay_incr;
elsif nramp = '0' and StoredData = "011010110111" then SHout <= '1' after delay1 + 1719*delay_incr;
elsif nramp = '0' and StoredData = "011010111000" then SHout <= '1' after delay1 + 1720*delay_incr;
elsif nramp = '0' and StoredData = "011010111001" then SHout <= '1' after delay1 + 1721*delay_incr;
elsif nramp = '0' and StoredData = "011010111010" then SHout <= '1' after delay1 + 1722*delay_incr;
elsif nramp = '0' and StoredData = "011010111011" then SHout <= '1' after delay1 + 1723*delay_incr;
elsif nramp = '0' and StoredData = "011010111100" then SHout <= '1' after delay1 + 1724*delay_incr;
elsif nramp = '0' and StoredData = "011010111101" then SHout <= '1' after delay1 + 1725*delay_incr;
elsif nramp = '0' and StoredData = "011010111110" then SHout <= '1' after delay1 + 1726*delay_incr;
elsif nramp = '0' and StoredData = "011010111111" then SHout <= '1' after delay1 + 1727*delay_incr;
elsif nramp = '0' and StoredData = "011011000000" then SHout <= '1' after delay1 + 1728*delay_incr;
elsif nramp = '0' and StoredData = "011011000001" then SHout <= '1' after delay1 + 1729*delay_incr;
elsif nramp = '0' and StoredData = "011011000010" then SHout <= '1' after delay1 + 1730*delay_incr;
elsif nramp = '0' and StoredData = "011011000011" then SHout <= '1' after delay1 + 1731*delay_incr;
elsif nramp = '0' and StoredData = "011011000100" then SHout <= '1' after delay1 + 1732*delay_incr;
elsif nramp = '0' and StoredData = "011011000101" then SHout <= '1' after delay1 + 1733*delay_incr;
elsif nramp = '0' and StoredData = "011011000110" then SHout <= '1' after delay1 + 1734*delay_incr;
elsif nramp = '0' and StoredData = "011011000111" then SHout <= '1' after delay1 + 1735*delay_incr;
elsif nramp = '0' and StoredData = "011011001000" then SHout <= '1' after delay1 + 1736*delay_incr;
elsif nramp = '0' and StoredData = "011011001001" then SHout <= '1' after delay1 + 1737*delay_incr;
elsif nramp = '0' and StoredData = "011011001010" then SHout <= '1' after delay1 + 1738*delay_incr;
elsif nramp = '0' and StoredData = "011011001011" then SHout <= '1' after delay1 + 1739*delay_incr;
elsif nramp = '0' and StoredData = "011011001100" then SHout <= '1' after delay1 + 1740*delay_incr;
elsif nramp = '0' and StoredData = "011011001101" then SHout <= '1' after delay1 + 1741*delay_incr;
elsif nramp = '0' and StoredData = "011011001110" then SHout <= '1' after delay1 + 1742*delay_incr;
elsif nramp = '0' and StoredData = "011011001111" then SHout <= '1' after delay1 + 1743*delay_incr;
elsif nramp = '0' and StoredData = "011011010000" then SHout <= '1' after delay1 + 1744*delay_incr;
elsif nramp = '0' and StoredData = "011011010001" then SHout <= '1' after delay1 + 1745*delay_incr;
elsif nramp = '0' and StoredData = "011011010010" then SHout <= '1' after delay1 + 1746*delay_incr;
elsif nramp = '0' and StoredData = "011011010011" then SHout <= '1' after delay1 + 1747*delay_incr;
elsif nramp = '0' and StoredData = "011011010100" then SHout <= '1' after delay1 + 1748*delay_incr;
elsif nramp = '0' and StoredData = "011011010101" then SHout <= '1' after delay1 + 1749*delay_incr;
elsif nramp = '0' and StoredData = "011011010110" then SHout <= '1' after delay1 + 1750*delay_incr;
elsif nramp = '0' and StoredData = "011011010111" then SHout <= '1' after delay1 + 1751*delay_incr;
elsif nramp = '0' and StoredData = "011011011000" then SHout <= '1' after delay1 + 1752*delay_incr;
elsif nramp = '0' and StoredData = "011011011001" then SHout <= '1' after delay1 + 1753*delay_incr;
elsif nramp = '0' and StoredData = "011011011010" then SHout <= '1' after delay1 + 1754*delay_incr;
elsif nramp = '0' and StoredData = "011011011011" then SHout <= '1' after delay1 + 1755*delay_incr;
elsif nramp = '0' and StoredData = "011011011100" then SHout <= '1' after delay1 + 1756*delay_incr;
elsif nramp = '0' and StoredData = "011011011101" then SHout <= '1' after delay1 + 1757*delay_incr;
elsif nramp = '0' and StoredData = "011011011110" then SHout <= '1' after delay1 + 1758*delay_incr;
elsif nramp = '0' and StoredData = "011011011111" then SHout <= '1' after delay1 + 1759*delay_incr;
elsif nramp = '0' and StoredData = "011011100000" then SHout <= '1' after delay1 + 1760*delay_incr;
elsif nramp = '0' and StoredData = "011011100001" then SHout <= '1' after delay1 + 1761*delay_incr;
elsif nramp = '0' and StoredData = "011011100010" then SHout <= '1' after delay1 + 1762*delay_incr;
elsif nramp = '0' and StoredData = "011011100011" then SHout <= '1' after delay1 + 1763*delay_incr;
elsif nramp = '0' and StoredData = "011011100100" then SHout <= '1' after delay1 + 1764*delay_incr;
elsif nramp = '0' and StoredData = "011011100101" then SHout <= '1' after delay1 + 1765*delay_incr;
elsif nramp = '0' and StoredData = "011011100110" then SHout <= '1' after delay1 + 1766*delay_incr;
elsif nramp = '0' and StoredData = "011011100111" then SHout <= '1' after delay1 + 1767*delay_incr;
elsif nramp = '0' and StoredData = "011011101000" then SHout <= '1' after delay1 + 1768*delay_incr;
elsif nramp = '0' and StoredData = "011011101001" then SHout <= '1' after delay1 + 1769*delay_incr;
elsif nramp = '0' and StoredData = "011011101010" then SHout <= '1' after delay1 + 1770*delay_incr;
elsif nramp = '0' and StoredData = "011011101011" then SHout <= '1' after delay1 + 1771*delay_incr;
elsif nramp = '0' and StoredData = "011011101100" then SHout <= '1' after delay1 + 1772*delay_incr;
elsif nramp = '0' and StoredData = "011011101101" then SHout <= '1' after delay1 + 1773*delay_incr;
elsif nramp = '0' and StoredData = "011011101110" then SHout <= '1' after delay1 + 1774*delay_incr;
elsif nramp = '0' and StoredData = "011011101111" then SHout <= '1' after delay1 + 1775*delay_incr;
elsif nramp = '0' and StoredData = "011011110000" then SHout <= '1' after delay1 + 1776*delay_incr;
elsif nramp = '0' and StoredData = "011011110001" then SHout <= '1' after delay1 + 1777*delay_incr;
elsif nramp = '0' and StoredData = "011011110010" then SHout <= '1' after delay1 + 1778*delay_incr;
elsif nramp = '0' and StoredData = "011011110011" then SHout <= '1' after delay1 + 1779*delay_incr;
elsif nramp = '0' and StoredData = "011011110100" then SHout <= '1' after delay1 + 1780*delay_incr;
elsif nramp = '0' and StoredData = "011011110101" then SHout <= '1' after delay1 + 1781*delay_incr;
elsif nramp = '0' and StoredData = "011011110110" then SHout <= '1' after delay1 + 1782*delay_incr;
elsif nramp = '0' and StoredData = "011011110111" then SHout <= '1' after delay1 + 1783*delay_incr;
elsif nramp = '0' and StoredData = "011011111000" then SHout <= '1' after delay1 + 1784*delay_incr;
elsif nramp = '0' and StoredData = "011011111001" then SHout <= '1' after delay1 + 1785*delay_incr;
elsif nramp = '0' and StoredData = "011011111010" then SHout <= '1' after delay1 + 1786*delay_incr;
elsif nramp = '0' and StoredData = "011011111011" then SHout <= '1' after delay1 + 1787*delay_incr;
elsif nramp = '0' and StoredData = "011011111100" then SHout <= '1' after delay1 + 1788*delay_incr;
elsif nramp = '0' and StoredData = "011011111101" then SHout <= '1' after delay1 + 1789*delay_incr;
elsif nramp = '0' and StoredData = "011011111110" then SHout <= '1' after delay1 + 1790*delay_incr;
elsif nramp = '0' and StoredData = "011011111111" then SHout <= '1' after delay1 + 1791*delay_incr;
elsif nramp = '0' and StoredData = "011100000000" then SHout <= '1' after delay1 + 1792*delay_incr;
elsif nramp = '0' and StoredData = "011100000001" then SHout <= '1' after delay1 + 1793*delay_incr;
elsif nramp = '0' and StoredData = "011100000010" then SHout <= '1' after delay1 + 1794*delay_incr;
elsif nramp = '0' and StoredData = "011100000011" then SHout <= '1' after delay1 + 1795*delay_incr;
elsif nramp = '0' and StoredData = "011100000100" then SHout <= '1' after delay1 + 1796*delay_incr;
elsif nramp = '0' and StoredData = "011100000101" then SHout <= '1' after delay1 + 1797*delay_incr;
elsif nramp = '0' and StoredData = "011100000110" then SHout <= '1' after delay1 + 1798*delay_incr;
elsif nramp = '0' and StoredData = "011100000111" then SHout <= '1' after delay1 + 1799*delay_incr;
elsif nramp = '0' and StoredData = "011100001000" then SHout <= '1' after delay1 + 1800*delay_incr;
elsif nramp = '0' and StoredData = "011100001001" then SHout <= '1' after delay1 + 1801*delay_incr;
elsif nramp = '0' and StoredData = "011100001010" then SHout <= '1' after delay1 + 1802*delay_incr;
elsif nramp = '0' and StoredData = "011100001011" then SHout <= '1' after delay1 + 1803*delay_incr;
elsif nramp = '0' and StoredData = "011100001100" then SHout <= '1' after delay1 + 1804*delay_incr;
elsif nramp = '0' and StoredData = "011100001101" then SHout <= '1' after delay1 + 1805*delay_incr;
elsif nramp = '0' and StoredData = "011100001110" then SHout <= '1' after delay1 + 1806*delay_incr;
elsif nramp = '0' and StoredData = "011100001111" then SHout <= '1' after delay1 + 1807*delay_incr;
elsif nramp = '0' and StoredData = "011100010000" then SHout <= '1' after delay1 + 1808*delay_incr;
elsif nramp = '0' and StoredData = "011100010001" then SHout <= '1' after delay1 + 1809*delay_incr;
elsif nramp = '0' and StoredData = "011100010010" then SHout <= '1' after delay1 + 1810*delay_incr;
elsif nramp = '0' and StoredData = "011100010011" then SHout <= '1' after delay1 + 1811*delay_incr;
elsif nramp = '0' and StoredData = "011100010100" then SHout <= '1' after delay1 + 1812*delay_incr;
elsif nramp = '0' and StoredData = "011100010101" then SHout <= '1' after delay1 + 1813*delay_incr;
elsif nramp = '0' and StoredData = "011100010110" then SHout <= '1' after delay1 + 1814*delay_incr;
elsif nramp = '0' and StoredData = "011100010111" then SHout <= '1' after delay1 + 1815*delay_incr;
elsif nramp = '0' and StoredData = "011100011000" then SHout <= '1' after delay1 + 1816*delay_incr;
elsif nramp = '0' and StoredData = "011100011001" then SHout <= '1' after delay1 + 1817*delay_incr;
elsif nramp = '0' and StoredData = "011100011010" then SHout <= '1' after delay1 + 1818*delay_incr;
elsif nramp = '0' and StoredData = "011100011011" then SHout <= '1' after delay1 + 1819*delay_incr;
elsif nramp = '0' and StoredData = "011100011100" then SHout <= '1' after delay1 + 1820*delay_incr;
elsif nramp = '0' and StoredData = "011100011101" then SHout <= '1' after delay1 + 1821*delay_incr;
elsif nramp = '0' and StoredData = "011100011110" then SHout <= '1' after delay1 + 1822*delay_incr;
elsif nramp = '0' and StoredData = "011100011111" then SHout <= '1' after delay1 + 1823*delay_incr;
elsif nramp = '0' and StoredData = "011100100000" then SHout <= '1' after delay1 + 1824*delay_incr;
elsif nramp = '0' and StoredData = "011100100001" then SHout <= '1' after delay1 + 1825*delay_incr;
elsif nramp = '0' and StoredData = "011100100010" then SHout <= '1' after delay1 + 1826*delay_incr;
elsif nramp = '0' and StoredData = "011100100011" then SHout <= '1' after delay1 + 1827*delay_incr;
elsif nramp = '0' and StoredData = "011100100100" then SHout <= '1' after delay1 + 1828*delay_incr;
elsif nramp = '0' and StoredData = "011100100101" then SHout <= '1' after delay1 + 1829*delay_incr;
elsif nramp = '0' and StoredData = "011100100110" then SHout <= '1' after delay1 + 1830*delay_incr;
elsif nramp = '0' and StoredData = "011100100111" then SHout <= '1' after delay1 + 1831*delay_incr;
elsif nramp = '0' and StoredData = "011100101000" then SHout <= '1' after delay1 + 1832*delay_incr;
elsif nramp = '0' and StoredData = "011100101001" then SHout <= '1' after delay1 + 1833*delay_incr;
elsif nramp = '0' and StoredData = "011100101010" then SHout <= '1' after delay1 + 1834*delay_incr;
elsif nramp = '0' and StoredData = "011100101011" then SHout <= '1' after delay1 + 1835*delay_incr;
elsif nramp = '0' and StoredData = "011100101100" then SHout <= '1' after delay1 + 1836*delay_incr;
elsif nramp = '0' and StoredData = "011100101101" then SHout <= '1' after delay1 + 1837*delay_incr;
elsif nramp = '0' and StoredData = "011100101110" then SHout <= '1' after delay1 + 1838*delay_incr;
elsif nramp = '0' and StoredData = "011100101111" then SHout <= '1' after delay1 + 1839*delay_incr;
elsif nramp = '0' and StoredData = "011100110000" then SHout <= '1' after delay1 + 1840*delay_incr;
elsif nramp = '0' and StoredData = "011100110001" then SHout <= '1' after delay1 + 1841*delay_incr;
elsif nramp = '0' and StoredData = "011100110010" then SHout <= '1' after delay1 + 1842*delay_incr;
elsif nramp = '0' and StoredData = "011100110011" then SHout <= '1' after delay1 + 1843*delay_incr;
elsif nramp = '0' and StoredData = "011100110100" then SHout <= '1' after delay1 + 1844*delay_incr;
elsif nramp = '0' and StoredData = "011100110101" then SHout <= '1' after delay1 + 1845*delay_incr;
elsif nramp = '0' and StoredData = "011100110110" then SHout <= '1' after delay1 + 1846*delay_incr;
elsif nramp = '0' and StoredData = "011100110111" then SHout <= '1' after delay1 + 1847*delay_incr;
elsif nramp = '0' and StoredData = "011100111000" then SHout <= '1' after delay1 + 1848*delay_incr;
elsif nramp = '0' and StoredData = "011100111001" then SHout <= '1' after delay1 + 1849*delay_incr;
elsif nramp = '0' and StoredData = "011100111010" then SHout <= '1' after delay1 + 1850*delay_incr;
elsif nramp = '0' and StoredData = "011100111011" then SHout <= '1' after delay1 + 1851*delay_incr;
elsif nramp = '0' and StoredData = "011100111100" then SHout <= '1' after delay1 + 1852*delay_incr;
elsif nramp = '0' and StoredData = "011100111101" then SHout <= '1' after delay1 + 1853*delay_incr;
elsif nramp = '0' and StoredData = "011100111110" then SHout <= '1' after delay1 + 1854*delay_incr;
elsif nramp = '0' and StoredData = "011100111111" then SHout <= '1' after delay1 + 1855*delay_incr;
elsif nramp = '0' and StoredData = "011101000000" then SHout <= '1' after delay1 + 1856*delay_incr;
elsif nramp = '0' and StoredData = "011101000001" then SHout <= '1' after delay1 + 1857*delay_incr;
elsif nramp = '0' and StoredData = "011101000010" then SHout <= '1' after delay1 + 1858*delay_incr;
elsif nramp = '0' and StoredData = "011101000011" then SHout <= '1' after delay1 + 1859*delay_incr;
elsif nramp = '0' and StoredData = "011101000100" then SHout <= '1' after delay1 + 1860*delay_incr;
elsif nramp = '0' and StoredData = "011101000101" then SHout <= '1' after delay1 + 1861*delay_incr;
elsif nramp = '0' and StoredData = "011101000110" then SHout <= '1' after delay1 + 1862*delay_incr;
elsif nramp = '0' and StoredData = "011101000111" then SHout <= '1' after delay1 + 1863*delay_incr;
elsif nramp = '0' and StoredData = "011101001000" then SHout <= '1' after delay1 + 1864*delay_incr;
elsif nramp = '0' and StoredData = "011101001001" then SHout <= '1' after delay1 + 1865*delay_incr;
elsif nramp = '0' and StoredData = "011101001010" then SHout <= '1' after delay1 + 1866*delay_incr;
elsif nramp = '0' and StoredData = "011101001011" then SHout <= '1' after delay1 + 1867*delay_incr;
elsif nramp = '0' and StoredData = "011101001100" then SHout <= '1' after delay1 + 1868*delay_incr;
elsif nramp = '0' and StoredData = "011101001101" then SHout <= '1' after delay1 + 1869*delay_incr;
elsif nramp = '0' and StoredData = "011101001110" then SHout <= '1' after delay1 + 1870*delay_incr;
elsif nramp = '0' and StoredData = "011101001111" then SHout <= '1' after delay1 + 1871*delay_incr;
elsif nramp = '0' and StoredData = "011101010000" then SHout <= '1' after delay1 + 1872*delay_incr;
elsif nramp = '0' and StoredData = "011101010001" then SHout <= '1' after delay1 + 1873*delay_incr;
elsif nramp = '0' and StoredData = "011101010010" then SHout <= '1' after delay1 + 1874*delay_incr;
elsif nramp = '0' and StoredData = "011101010011" then SHout <= '1' after delay1 + 1875*delay_incr;
elsif nramp = '0' and StoredData = "011101010100" then SHout <= '1' after delay1 + 1876*delay_incr;
elsif nramp = '0' and StoredData = "011101010101" then SHout <= '1' after delay1 + 1877*delay_incr;
elsif nramp = '0' and StoredData = "011101010110" then SHout <= '1' after delay1 + 1878*delay_incr;
elsif nramp = '0' and StoredData = "011101010111" then SHout <= '1' after delay1 + 1879*delay_incr;
elsif nramp = '0' and StoredData = "011101011000" then SHout <= '1' after delay1 + 1880*delay_incr;
elsif nramp = '0' and StoredData = "011101011001" then SHout <= '1' after delay1 + 1881*delay_incr;
elsif nramp = '0' and StoredData = "011101011010" then SHout <= '1' after delay1 + 1882*delay_incr;
elsif nramp = '0' and StoredData = "011101011011" then SHout <= '1' after delay1 + 1883*delay_incr;
elsif nramp = '0' and StoredData = "011101011100" then SHout <= '1' after delay1 + 1884*delay_incr;
elsif nramp = '0' and StoredData = "011101011101" then SHout <= '1' after delay1 + 1885*delay_incr;
elsif nramp = '0' and StoredData = "011101011110" then SHout <= '1' after delay1 + 1886*delay_incr;
elsif nramp = '0' and StoredData = "011101011111" then SHout <= '1' after delay1 + 1887*delay_incr;
elsif nramp = '0' and StoredData = "011101100000" then SHout <= '1' after delay1 + 1888*delay_incr;
elsif nramp = '0' and StoredData = "011101100001" then SHout <= '1' after delay1 + 1889*delay_incr;
elsif nramp = '0' and StoredData = "011101100010" then SHout <= '1' after delay1 + 1890*delay_incr;
elsif nramp = '0' and StoredData = "011101100011" then SHout <= '1' after delay1 + 1891*delay_incr;
elsif nramp = '0' and StoredData = "011101100100" then SHout <= '1' after delay1 + 1892*delay_incr;
elsif nramp = '0' and StoredData = "011101100101" then SHout <= '1' after delay1 + 1893*delay_incr;
elsif nramp = '0' and StoredData = "011101100110" then SHout <= '1' after delay1 + 1894*delay_incr;
elsif nramp = '0' and StoredData = "011101100111" then SHout <= '1' after delay1 + 1895*delay_incr;
elsif nramp = '0' and StoredData = "011101101000" then SHout <= '1' after delay1 + 1896*delay_incr;
elsif nramp = '0' and StoredData = "011101101001" then SHout <= '1' after delay1 + 1897*delay_incr;
elsif nramp = '0' and StoredData = "011101101010" then SHout <= '1' after delay1 + 1898*delay_incr;
elsif nramp = '0' and StoredData = "011101101011" then SHout <= '1' after delay1 + 1899*delay_incr;
elsif nramp = '0' and StoredData = "011101101100" then SHout <= '1' after delay1 + 1900*delay_incr;
elsif nramp = '0' and StoredData = "011101101101" then SHout <= '1' after delay1 + 1901*delay_incr;
elsif nramp = '0' and StoredData = "011101101110" then SHout <= '1' after delay1 + 1902*delay_incr;
elsif nramp = '0' and StoredData = "011101101111" then SHout <= '1' after delay1 + 1903*delay_incr;
elsif nramp = '0' and StoredData = "011101110000" then SHout <= '1' after delay1 + 1904*delay_incr;
elsif nramp = '0' and StoredData = "011101110001" then SHout <= '1' after delay1 + 1905*delay_incr;
elsif nramp = '0' and StoredData = "011101110010" then SHout <= '1' after delay1 + 1906*delay_incr;
elsif nramp = '0' and StoredData = "011101110011" then SHout <= '1' after delay1 + 1907*delay_incr;
elsif nramp = '0' and StoredData = "011101110100" then SHout <= '1' after delay1 + 1908*delay_incr;
elsif nramp = '0' and StoredData = "011101110101" then SHout <= '1' after delay1 + 1909*delay_incr;
elsif nramp = '0' and StoredData = "011101110110" then SHout <= '1' after delay1 + 1910*delay_incr;
elsif nramp = '0' and StoredData = "011101110111" then SHout <= '1' after delay1 + 1911*delay_incr;
elsif nramp = '0' and StoredData = "011101111000" then SHout <= '1' after delay1 + 1912*delay_incr;
elsif nramp = '0' and StoredData = "011101111001" then SHout <= '1' after delay1 + 1913*delay_incr;
elsif nramp = '0' and StoredData = "011101111010" then SHout <= '1' after delay1 + 1914*delay_incr;
elsif nramp = '0' and StoredData = "011101111011" then SHout <= '1' after delay1 + 1915*delay_incr;
elsif nramp = '0' and StoredData = "011101111100" then SHout <= '1' after delay1 + 1916*delay_incr;
elsif nramp = '0' and StoredData = "011101111101" then SHout <= '1' after delay1 + 1917*delay_incr;
elsif nramp = '0' and StoredData = "011101111110" then SHout <= '1' after delay1 + 1918*delay_incr;
elsif nramp = '0' and StoredData = "011101111111" then SHout <= '1' after delay1 + 1919*delay_incr;
elsif nramp = '0' and StoredData = "011110000000" then SHout <= '1' after delay1 + 1920*delay_incr;
elsif nramp = '0' and StoredData = "011110000001" then SHout <= '1' after delay1 + 1921*delay_incr;
elsif nramp = '0' and StoredData = "011110000010" then SHout <= '1' after delay1 + 1922*delay_incr;
elsif nramp = '0' and StoredData = "011110000011" then SHout <= '1' after delay1 + 1923*delay_incr;
elsif nramp = '0' and StoredData = "011110000100" then SHout <= '1' after delay1 + 1924*delay_incr;
elsif nramp = '0' and StoredData = "011110000101" then SHout <= '1' after delay1 + 1925*delay_incr;
elsif nramp = '0' and StoredData = "011110000110" then SHout <= '1' after delay1 + 1926*delay_incr;
elsif nramp = '0' and StoredData = "011110000111" then SHout <= '1' after delay1 + 1927*delay_incr;
elsif nramp = '0' and StoredData = "011110001000" then SHout <= '1' after delay1 + 1928*delay_incr;
elsif nramp = '0' and StoredData = "011110001001" then SHout <= '1' after delay1 + 1929*delay_incr;
elsif nramp = '0' and StoredData = "011110001010" then SHout <= '1' after delay1 + 1930*delay_incr;
elsif nramp = '0' and StoredData = "011110001011" then SHout <= '1' after delay1 + 1931*delay_incr;
elsif nramp = '0' and StoredData = "011110001100" then SHout <= '1' after delay1 + 1932*delay_incr;
elsif nramp = '0' and StoredData = "011110001101" then SHout <= '1' after delay1 + 1933*delay_incr;
elsif nramp = '0' and StoredData = "011110001110" then SHout <= '1' after delay1 + 1934*delay_incr;
elsif nramp = '0' and StoredData = "011110001111" then SHout <= '1' after delay1 + 1935*delay_incr;
elsif nramp = '0' and StoredData = "011110010000" then SHout <= '1' after delay1 + 1936*delay_incr;
elsif nramp = '0' and StoredData = "011110010001" then SHout <= '1' after delay1 + 1937*delay_incr;
elsif nramp = '0' and StoredData = "011110010010" then SHout <= '1' after delay1 + 1938*delay_incr;
elsif nramp = '0' and StoredData = "011110010011" then SHout <= '1' after delay1 + 1939*delay_incr;
elsif nramp = '0' and StoredData = "011110010100" then SHout <= '1' after delay1 + 1940*delay_incr;
elsif nramp = '0' and StoredData = "011110010101" then SHout <= '1' after delay1 + 1941*delay_incr;
elsif nramp = '0' and StoredData = "011110010110" then SHout <= '1' after delay1 + 1942*delay_incr;
elsif nramp = '0' and StoredData = "011110010111" then SHout <= '1' after delay1 + 1943*delay_incr;
elsif nramp = '0' and StoredData = "011110011000" then SHout <= '1' after delay1 + 1944*delay_incr;
elsif nramp = '0' and StoredData = "011110011001" then SHout <= '1' after delay1 + 1945*delay_incr;
elsif nramp = '0' and StoredData = "011110011010" then SHout <= '1' after delay1 + 1946*delay_incr;
elsif nramp = '0' and StoredData = "011110011011" then SHout <= '1' after delay1 + 1947*delay_incr;
elsif nramp = '0' and StoredData = "011110011100" then SHout <= '1' after delay1 + 1948*delay_incr;
elsif nramp = '0' and StoredData = "011110011101" then SHout <= '1' after delay1 + 1949*delay_incr;
elsif nramp = '0' and StoredData = "011110011110" then SHout <= '1' after delay1 + 1950*delay_incr;
elsif nramp = '0' and StoredData = "011110011111" then SHout <= '1' after delay1 + 1951*delay_incr;
elsif nramp = '0' and StoredData = "011110100000" then SHout <= '1' after delay1 + 1952*delay_incr;
elsif nramp = '0' and StoredData = "011110100001" then SHout <= '1' after delay1 + 1953*delay_incr;
elsif nramp = '0' and StoredData = "011110100010" then SHout <= '1' after delay1 + 1954*delay_incr;
elsif nramp = '0' and StoredData = "011110100011" then SHout <= '1' after delay1 + 1955*delay_incr;
elsif nramp = '0' and StoredData = "011110100100" then SHout <= '1' after delay1 + 1956*delay_incr;
elsif nramp = '0' and StoredData = "011110100101" then SHout <= '1' after delay1 + 1957*delay_incr;
elsif nramp = '0' and StoredData = "011110100110" then SHout <= '1' after delay1 + 1958*delay_incr;
elsif nramp = '0' and StoredData = "011110100111" then SHout <= '1' after delay1 + 1959*delay_incr;
elsif nramp = '0' and StoredData = "011110101000" then SHout <= '1' after delay1 + 1960*delay_incr;
elsif nramp = '0' and StoredData = "011110101001" then SHout <= '1' after delay1 + 1961*delay_incr;
elsif nramp = '0' and StoredData = "011110101010" then SHout <= '1' after delay1 + 1962*delay_incr;
elsif nramp = '0' and StoredData = "011110101011" then SHout <= '1' after delay1 + 1963*delay_incr;
elsif nramp = '0' and StoredData = "011110101100" then SHout <= '1' after delay1 + 1964*delay_incr;
elsif nramp = '0' and StoredData = "011110101101" then SHout <= '1' after delay1 + 1965*delay_incr;
elsif nramp = '0' and StoredData = "011110101110" then SHout <= '1' after delay1 + 1966*delay_incr;
elsif nramp = '0' and StoredData = "011110101111" then SHout <= '1' after delay1 + 1967*delay_incr;
elsif nramp = '0' and StoredData = "011110110000" then SHout <= '1' after delay1 + 1968*delay_incr;
elsif nramp = '0' and StoredData = "011110110001" then SHout <= '1' after delay1 + 1969*delay_incr;
elsif nramp = '0' and StoredData = "011110110010" then SHout <= '1' after delay1 + 1970*delay_incr;
elsif nramp = '0' and StoredData = "011110110011" then SHout <= '1' after delay1 + 1971*delay_incr;
elsif nramp = '0' and StoredData = "011110110100" then SHout <= '1' after delay1 + 1972*delay_incr;
elsif nramp = '0' and StoredData = "011110110101" then SHout <= '1' after delay1 + 1973*delay_incr;
elsif nramp = '0' and StoredData = "011110110110" then SHout <= '1' after delay1 + 1974*delay_incr;
elsif nramp = '0' and StoredData = "011110110111" then SHout <= '1' after delay1 + 1975*delay_incr;
elsif nramp = '0' and StoredData = "011110111000" then SHout <= '1' after delay1 + 1976*delay_incr;
elsif nramp = '0' and StoredData = "011110111001" then SHout <= '1' after delay1 + 1977*delay_incr;
elsif nramp = '0' and StoredData = "011110111010" then SHout <= '1' after delay1 + 1978*delay_incr;
elsif nramp = '0' and StoredData = "011110111011" then SHout <= '1' after delay1 + 1979*delay_incr;
elsif nramp = '0' and StoredData = "011110111100" then SHout <= '1' after delay1 + 1980*delay_incr;
elsif nramp = '0' and StoredData = "011110111101" then SHout <= '1' after delay1 + 1981*delay_incr;
elsif nramp = '0' and StoredData = "011110111110" then SHout <= '1' after delay1 + 1982*delay_incr;
elsif nramp = '0' and StoredData = "011110111111" then SHout <= '1' after delay1 + 1983*delay_incr;
elsif nramp = '0' and StoredData = "011111000000" then SHout <= '1' after delay1 + 1984*delay_incr;
elsif nramp = '0' and StoredData = "011111000001" then SHout <= '1' after delay1 + 1985*delay_incr;
elsif nramp = '0' and StoredData = "011111000010" then SHout <= '1' after delay1 + 1986*delay_incr;
elsif nramp = '0' and StoredData = "011111000011" then SHout <= '1' after delay1 + 1987*delay_incr;
elsif nramp = '0' and StoredData = "011111000100" then SHout <= '1' after delay1 + 1988*delay_incr;
elsif nramp = '0' and StoredData = "011111000101" then SHout <= '1' after delay1 + 1989*delay_incr;
elsif nramp = '0' and StoredData = "011111000110" then SHout <= '1' after delay1 + 1990*delay_incr;
elsif nramp = '0' and StoredData = "011111000111" then SHout <= '1' after delay1 + 1991*delay_incr;
elsif nramp = '0' and StoredData = "011111001000" then SHout <= '1' after delay1 + 1992*delay_incr;
elsif nramp = '0' and StoredData = "011111001001" then SHout <= '1' after delay1 + 1993*delay_incr;
elsif nramp = '0' and StoredData = "011111001010" then SHout <= '1' after delay1 + 1994*delay_incr;
elsif nramp = '0' and StoredData = "011111001011" then SHout <= '1' after delay1 + 1995*delay_incr;
elsif nramp = '0' and StoredData = "011111001100" then SHout <= '1' after delay1 + 1996*delay_incr;
elsif nramp = '0' and StoredData = "011111001101" then SHout <= '1' after delay1 + 1997*delay_incr;
elsif nramp = '0' and StoredData = "011111001110" then SHout <= '1' after delay1 + 1998*delay_incr;
elsif nramp = '0' and StoredData = "011111001111" then SHout <= '1' after delay1 + 1999*delay_incr;
elsif nramp = '0' and StoredData = "011111010000" then SHout <= '1' after delay1 + 2000*delay_incr;
elsif nramp = '0' and StoredData = "011111010001" then SHout <= '1' after delay1 + 2001*delay_incr;
elsif nramp = '0' and StoredData = "011111010010" then SHout <= '1' after delay1 + 2002*delay_incr;
elsif nramp = '0' and StoredData = "011111010011" then SHout <= '1' after delay1 + 2003*delay_incr;
elsif nramp = '0' and StoredData = "011111010100" then SHout <= '1' after delay1 + 2004*delay_incr;
elsif nramp = '0' and StoredData = "011111010101" then SHout <= '1' after delay1 + 2005*delay_incr;
elsif nramp = '0' and StoredData = "011111010110" then SHout <= '1' after delay1 + 2006*delay_incr;
elsif nramp = '0' and StoredData = "011111010111" then SHout <= '1' after delay1 + 2007*delay_incr;
elsif nramp = '0' and StoredData = "011111011000" then SHout <= '1' after delay1 + 2008*delay_incr;
elsif nramp = '0' and StoredData = "011111011001" then SHout <= '1' after delay1 + 2009*delay_incr;
elsif nramp = '0' and StoredData = "011111011010" then SHout <= '1' after delay1 + 2010*delay_incr;
elsif nramp = '0' and StoredData = "011111011011" then SHout <= '1' after delay1 + 2011*delay_incr;
elsif nramp = '0' and StoredData = "011111011100" then SHout <= '1' after delay1 + 2012*delay_incr;
elsif nramp = '0' and StoredData = "011111011101" then SHout <= '1' after delay1 + 2013*delay_incr;
elsif nramp = '0' and StoredData = "011111011110" then SHout <= '1' after delay1 + 2014*delay_incr;
elsif nramp = '0' and StoredData = "011111011111" then SHout <= '1' after delay1 + 2015*delay_incr;
elsif nramp = '0' and StoredData = "011111100000" then SHout <= '1' after delay1 + 2016*delay_incr;
elsif nramp = '0' and StoredData = "011111100001" then SHout <= '1' after delay1 + 2017*delay_incr;
elsif nramp = '0' and StoredData = "011111100010" then SHout <= '1' after delay1 + 2018*delay_incr;
elsif nramp = '0' and StoredData = "011111100011" then SHout <= '1' after delay1 + 2019*delay_incr;
elsif nramp = '0' and StoredData = "011111100100" then SHout <= '1' after delay1 + 2020*delay_incr;
elsif nramp = '0' and StoredData = "011111100101" then SHout <= '1' after delay1 + 2021*delay_incr;
elsif nramp = '0' and StoredData = "011111100110" then SHout <= '1' after delay1 + 2022*delay_incr;
elsif nramp = '0' and StoredData = "011111100111" then SHout <= '1' after delay1 + 2023*delay_incr;
elsif nramp = '0' and StoredData = "011111101000" then SHout <= '1' after delay1 + 2024*delay_incr;
elsif nramp = '0' and StoredData = "011111101001" then SHout <= '1' after delay1 + 2025*delay_incr;
elsif nramp = '0' and StoredData = "011111101010" then SHout <= '1' after delay1 + 2026*delay_incr;
elsif nramp = '0' and StoredData = "011111101011" then SHout <= '1' after delay1 + 2027*delay_incr;
elsif nramp = '0' and StoredData = "011111101100" then SHout <= '1' after delay1 + 2028*delay_incr;
elsif nramp = '0' and StoredData = "011111101101" then SHout <= '1' after delay1 + 2029*delay_incr;
elsif nramp = '0' and StoredData = "011111101110" then SHout <= '1' after delay1 + 2030*delay_incr;
elsif nramp = '0' and StoredData = "011111101111" then SHout <= '1' after delay1 + 2031*delay_incr;
elsif nramp = '0' and StoredData = "011111110000" then SHout <= '1' after delay1 + 2032*delay_incr;
elsif nramp = '0' and StoredData = "011111110001" then SHout <= '1' after delay1 + 2033*delay_incr;
elsif nramp = '0' and StoredData = "011111110010" then SHout <= '1' after delay1 + 2034*delay_incr;
elsif nramp = '0' and StoredData = "011111110011" then SHout <= '1' after delay1 + 2035*delay_incr;
elsif nramp = '0' and StoredData = "011111110100" then SHout <= '1' after delay1 + 2036*delay_incr;
elsif nramp = '0' and StoredData = "011111110101" then SHout <= '1' after delay1 + 2037*delay_incr;
elsif nramp = '0' and StoredData = "011111110110" then SHout <= '1' after delay1 + 2038*delay_incr;
elsif nramp = '0' and StoredData = "011111110111" then SHout <= '1' after delay1 + 2039*delay_incr;
elsif nramp = '0' and StoredData = "011111111000" then SHout <= '1' after delay1 + 2040*delay_incr;
elsif nramp = '0' and StoredData = "011111111001" then SHout <= '1' after delay1 + 2041*delay_incr;
elsif nramp = '0' and StoredData = "011111111010" then SHout <= '1' after delay1 + 2042*delay_incr;
elsif nramp = '0' and StoredData = "011111111011" then SHout <= '1' after delay1 + 2043*delay_incr;
elsif nramp = '0' and StoredData = "011111111100" then SHout <= '1' after delay1 + 2044*delay_incr;
elsif nramp = '0' and StoredData = "011111111101" then SHout <= '1' after delay1 + 2045*delay_incr;
elsif nramp = '0' and StoredData = "011111111110" then SHout <= '1' after delay1 + 2046*delay_incr;
elsif nramp = '0' and StoredData = "011111111111" then SHout <= '1' after delay1 + 2047*delay_incr;
elsif nramp = '0' and StoredData = "100000000000" then SHout <= '1' after delay1 + 2048*delay_incr;
elsif nramp = '0' and StoredData = "100000000001" then SHout <= '1' after delay1 + 2049*delay_incr;
elsif nramp = '0' and StoredData = "100000000010" then SHout <= '1' after delay1 + 2050*delay_incr;
elsif nramp = '0' and StoredData = "100000000011" then SHout <= '1' after delay1 + 2051*delay_incr;
elsif nramp = '0' and StoredData = "100000000100" then SHout <= '1' after delay1 + 2052*delay_incr;
elsif nramp = '0' and StoredData = "100000000101" then SHout <= '1' after delay1 + 2053*delay_incr;
elsif nramp = '0' and StoredData = "100000000110" then SHout <= '1' after delay1 + 2054*delay_incr;
elsif nramp = '0' and StoredData = "100000000111" then SHout <= '1' after delay1 + 2055*delay_incr;
elsif nramp = '0' and StoredData = "100000001000" then SHout <= '1' after delay1 + 2056*delay_incr;
elsif nramp = '0' and StoredData = "100000001001" then SHout <= '1' after delay1 + 2057*delay_incr;
elsif nramp = '0' and StoredData = "100000001010" then SHout <= '1' after delay1 + 2058*delay_incr;
elsif nramp = '0' and StoredData = "100000001011" then SHout <= '1' after delay1 + 2059*delay_incr;
elsif nramp = '0' and StoredData = "100000001100" then SHout <= '1' after delay1 + 2060*delay_incr;
elsif nramp = '0' and StoredData = "100000001101" then SHout <= '1' after delay1 + 2061*delay_incr;
elsif nramp = '0' and StoredData = "100000001110" then SHout <= '1' after delay1 + 2062*delay_incr;
elsif nramp = '0' and StoredData = "100000001111" then SHout <= '1' after delay1 + 2063*delay_incr;
elsif nramp = '0' and StoredData = "100000010000" then SHout <= '1' after delay1 + 2064*delay_incr;
elsif nramp = '0' and StoredData = "100000010001" then SHout <= '1' after delay1 + 2065*delay_incr;
elsif nramp = '0' and StoredData = "100000010010" then SHout <= '1' after delay1 + 2066*delay_incr;
elsif nramp = '0' and StoredData = "100000010011" then SHout <= '1' after delay1 + 2067*delay_incr;
elsif nramp = '0' and StoredData = "100000010100" then SHout <= '1' after delay1 + 2068*delay_incr;
elsif nramp = '0' and StoredData = "100000010101" then SHout <= '1' after delay1 + 2069*delay_incr;
elsif nramp = '0' and StoredData = "100000010110" then SHout <= '1' after delay1 + 2070*delay_incr;
elsif nramp = '0' and StoredData = "100000010111" then SHout <= '1' after delay1 + 2071*delay_incr;
elsif nramp = '0' and StoredData = "100000011000" then SHout <= '1' after delay1 + 2072*delay_incr;
elsif nramp = '0' and StoredData = "100000011001" then SHout <= '1' after delay1 + 2073*delay_incr;
elsif nramp = '0' and StoredData = "100000011010" then SHout <= '1' after delay1 + 2074*delay_incr;
elsif nramp = '0' and StoredData = "100000011011" then SHout <= '1' after delay1 + 2075*delay_incr;
elsif nramp = '0' and StoredData = "100000011100" then SHout <= '1' after delay1 + 2076*delay_incr;
elsif nramp = '0' and StoredData = "100000011101" then SHout <= '1' after delay1 + 2077*delay_incr;
elsif nramp = '0' and StoredData = "100000011110" then SHout <= '1' after delay1 + 2078*delay_incr;
elsif nramp = '0' and StoredData = "100000011111" then SHout <= '1' after delay1 + 2079*delay_incr;
elsif nramp = '0' and StoredData = "100000100000" then SHout <= '1' after delay1 + 2080*delay_incr;
elsif nramp = '0' and StoredData = "100000100001" then SHout <= '1' after delay1 + 2081*delay_incr;
elsif nramp = '0' and StoredData = "100000100010" then SHout <= '1' after delay1 + 2082*delay_incr;
elsif nramp = '0' and StoredData = "100000100011" then SHout <= '1' after delay1 + 2083*delay_incr;
elsif nramp = '0' and StoredData = "100000100100" then SHout <= '1' after delay1 + 2084*delay_incr;
elsif nramp = '0' and StoredData = "100000100101" then SHout <= '1' after delay1 + 2085*delay_incr;
elsif nramp = '0' and StoredData = "100000100110" then SHout <= '1' after delay1 + 2086*delay_incr;
elsif nramp = '0' and StoredData = "100000100111" then SHout <= '1' after delay1 + 2087*delay_incr;
elsif nramp = '0' and StoredData = "100000101000" then SHout <= '1' after delay1 + 2088*delay_incr;
elsif nramp = '0' and StoredData = "100000101001" then SHout <= '1' after delay1 + 2089*delay_incr;
elsif nramp = '0' and StoredData = "100000101010" then SHout <= '1' after delay1 + 2090*delay_incr;
elsif nramp = '0' and StoredData = "100000101011" then SHout <= '1' after delay1 + 2091*delay_incr;
elsif nramp = '0' and StoredData = "100000101100" then SHout <= '1' after delay1 + 2092*delay_incr;
elsif nramp = '0' and StoredData = "100000101101" then SHout <= '1' after delay1 + 2093*delay_incr;
elsif nramp = '0' and StoredData = "100000101110" then SHout <= '1' after delay1 + 2094*delay_incr;
elsif nramp = '0' and StoredData = "100000101111" then SHout <= '1' after delay1 + 2095*delay_incr;
elsif nramp = '0' and StoredData = "100000110000" then SHout <= '1' after delay1 + 2096*delay_incr;
elsif nramp = '0' and StoredData = "100000110001" then SHout <= '1' after delay1 + 2097*delay_incr;
elsif nramp = '0' and StoredData = "100000110010" then SHout <= '1' after delay1 + 2098*delay_incr;
elsif nramp = '0' and StoredData = "100000110011" then SHout <= '1' after delay1 + 2099*delay_incr;
elsif nramp = '0' and StoredData = "100000110100" then SHout <= '1' after delay1 + 2100*delay_incr;
elsif nramp = '0' and StoredData = "100000110101" then SHout <= '1' after delay1 + 2101*delay_incr;
elsif nramp = '0' and StoredData = "100000110110" then SHout <= '1' after delay1 + 2102*delay_incr;
elsif nramp = '0' and StoredData = "100000110111" then SHout <= '1' after delay1 + 2103*delay_incr;
elsif nramp = '0' and StoredData = "100000111000" then SHout <= '1' after delay1 + 2104*delay_incr;
elsif nramp = '0' and StoredData = "100000111001" then SHout <= '1' after delay1 + 2105*delay_incr;
elsif nramp = '0' and StoredData = "100000111010" then SHout <= '1' after delay1 + 2106*delay_incr;
elsif nramp = '0' and StoredData = "100000111011" then SHout <= '1' after delay1 + 2107*delay_incr;
elsif nramp = '0' and StoredData = "100000111100" then SHout <= '1' after delay1 + 2108*delay_incr;
elsif nramp = '0' and StoredData = "100000111101" then SHout <= '1' after delay1 + 2109*delay_incr;
elsif nramp = '0' and StoredData = "100000111110" then SHout <= '1' after delay1 + 2110*delay_incr;
elsif nramp = '0' and StoredData = "100000111111" then SHout <= '1' after delay1 + 2111*delay_incr;
elsif nramp = '0' and StoredData = "100001000000" then SHout <= '1' after delay1 + 2112*delay_incr;
elsif nramp = '0' and StoredData = "100001000001" then SHout <= '1' after delay1 + 2113*delay_incr;
elsif nramp = '0' and StoredData = "100001000010" then SHout <= '1' after delay1 + 2114*delay_incr;
elsif nramp = '0' and StoredData = "100001000011" then SHout <= '1' after delay1 + 2115*delay_incr;
elsif nramp = '0' and StoredData = "100001000100" then SHout <= '1' after delay1 + 2116*delay_incr;
elsif nramp = '0' and StoredData = "100001000101" then SHout <= '1' after delay1 + 2117*delay_incr;
elsif nramp = '0' and StoredData = "100001000110" then SHout <= '1' after delay1 + 2118*delay_incr;
elsif nramp = '0' and StoredData = "100001000111" then SHout <= '1' after delay1 + 2119*delay_incr;
elsif nramp = '0' and StoredData = "100001001000" then SHout <= '1' after delay1 + 2120*delay_incr;
elsif nramp = '0' and StoredData = "100001001001" then SHout <= '1' after delay1 + 2121*delay_incr;
elsif nramp = '0' and StoredData = "100001001010" then SHout <= '1' after delay1 + 2122*delay_incr;
elsif nramp = '0' and StoredData = "100001001011" then SHout <= '1' after delay1 + 2123*delay_incr;
elsif nramp = '0' and StoredData = "100001001100" then SHout <= '1' after delay1 + 2124*delay_incr;
elsif nramp = '0' and StoredData = "100001001101" then SHout <= '1' after delay1 + 2125*delay_incr;
elsif nramp = '0' and StoredData = "100001001110" then SHout <= '1' after delay1 + 2126*delay_incr;
elsif nramp = '0' and StoredData = "100001001111" then SHout <= '1' after delay1 + 2127*delay_incr;
elsif nramp = '0' and StoredData = "100001010000" then SHout <= '1' after delay1 + 2128*delay_incr;
elsif nramp = '0' and StoredData = "100001010001" then SHout <= '1' after delay1 + 2129*delay_incr;
elsif nramp = '0' and StoredData = "100001010010" then SHout <= '1' after delay1 + 2130*delay_incr;
elsif nramp = '0' and StoredData = "100001010011" then SHout <= '1' after delay1 + 2131*delay_incr;
elsif nramp = '0' and StoredData = "100001010100" then SHout <= '1' after delay1 + 2132*delay_incr;
elsif nramp = '0' and StoredData = "100001010101" then SHout <= '1' after delay1 + 2133*delay_incr;
elsif nramp = '0' and StoredData = "100001010110" then SHout <= '1' after delay1 + 2134*delay_incr;
elsif nramp = '0' and StoredData = "100001010111" then SHout <= '1' after delay1 + 2135*delay_incr;
elsif nramp = '0' and StoredData = "100001011000" then SHout <= '1' after delay1 + 2136*delay_incr;
elsif nramp = '0' and StoredData = "100001011001" then SHout <= '1' after delay1 + 2137*delay_incr;
elsif nramp = '0' and StoredData = "100001011010" then SHout <= '1' after delay1 + 2138*delay_incr;
elsif nramp = '0' and StoredData = "100001011011" then SHout <= '1' after delay1 + 2139*delay_incr;
elsif nramp = '0' and StoredData = "100001011100" then SHout <= '1' after delay1 + 2140*delay_incr;
elsif nramp = '0' and StoredData = "100001011101" then SHout <= '1' after delay1 + 2141*delay_incr;
elsif nramp = '0' and StoredData = "100001011110" then SHout <= '1' after delay1 + 2142*delay_incr;
elsif nramp = '0' and StoredData = "100001011111" then SHout <= '1' after delay1 + 2143*delay_incr;
elsif nramp = '0' and StoredData = "100001100000" then SHout <= '1' after delay1 + 2144*delay_incr;
elsif nramp = '0' and StoredData = "100001100001" then SHout <= '1' after delay1 + 2145*delay_incr;
elsif nramp = '0' and StoredData = "100001100010" then SHout <= '1' after delay1 + 2146*delay_incr;
elsif nramp = '0' and StoredData = "100001100011" then SHout <= '1' after delay1 + 2147*delay_incr;
elsif nramp = '0' and StoredData = "100001100100" then SHout <= '1' after delay1 + 2148*delay_incr;
elsif nramp = '0' and StoredData = "100001100101" then SHout <= '1' after delay1 + 2149*delay_incr;
elsif nramp = '0' and StoredData = "100001100110" then SHout <= '1' after delay1 + 2150*delay_incr;
elsif nramp = '0' and StoredData = "100001100111" then SHout <= '1' after delay1 + 2151*delay_incr;
elsif nramp = '0' and StoredData = "100001101000" then SHout <= '1' after delay1 + 2152*delay_incr;
elsif nramp = '0' and StoredData = "100001101001" then SHout <= '1' after delay1 + 2153*delay_incr;
elsif nramp = '0' and StoredData = "100001101010" then SHout <= '1' after delay1 + 2154*delay_incr;
elsif nramp = '0' and StoredData = "100001101011" then SHout <= '1' after delay1 + 2155*delay_incr;
elsif nramp = '0' and StoredData = "100001101100" then SHout <= '1' after delay1 + 2156*delay_incr;
elsif nramp = '0' and StoredData = "100001101101" then SHout <= '1' after delay1 + 2157*delay_incr;
elsif nramp = '0' and StoredData = "100001101110" then SHout <= '1' after delay1 + 2158*delay_incr;
elsif nramp = '0' and StoredData = "100001101111" then SHout <= '1' after delay1 + 2159*delay_incr;
elsif nramp = '0' and StoredData = "100001110000" then SHout <= '1' after delay1 + 2160*delay_incr;
elsif nramp = '0' and StoredData = "100001110001" then SHout <= '1' after delay1 + 2161*delay_incr;
elsif nramp = '0' and StoredData = "100001110010" then SHout <= '1' after delay1 + 2162*delay_incr;
elsif nramp = '0' and StoredData = "100001110011" then SHout <= '1' after delay1 + 2163*delay_incr;
elsif nramp = '0' and StoredData = "100001110100" then SHout <= '1' after delay1 + 2164*delay_incr;
elsif nramp = '0' and StoredData = "100001110101" then SHout <= '1' after delay1 + 2165*delay_incr;
elsif nramp = '0' and StoredData = "100001110110" then SHout <= '1' after delay1 + 2166*delay_incr;
elsif nramp = '0' and StoredData = "100001110111" then SHout <= '1' after delay1 + 2167*delay_incr;
elsif nramp = '0' and StoredData = "100001111000" then SHout <= '1' after delay1 + 2168*delay_incr;
elsif nramp = '0' and StoredData = "100001111001" then SHout <= '1' after delay1 + 2169*delay_incr;
elsif nramp = '0' and StoredData = "100001111010" then SHout <= '1' after delay1 + 2170*delay_incr;
elsif nramp = '0' and StoredData = "100001111011" then SHout <= '1' after delay1 + 2171*delay_incr;
elsif nramp = '0' and StoredData = "100001111100" then SHout <= '1' after delay1 + 2172*delay_incr;
elsif nramp = '0' and StoredData = "100001111101" then SHout <= '1' after delay1 + 2173*delay_incr;
elsif nramp = '0' and StoredData = "100001111110" then SHout <= '1' after delay1 + 2174*delay_incr;
elsif nramp = '0' and StoredData = "100001111111" then SHout <= '1' after delay1 + 2175*delay_incr;
elsif nramp = '0' and StoredData = "100010000000" then SHout <= '1' after delay1 + 2176*delay_incr;
elsif nramp = '0' and StoredData = "100010000001" then SHout <= '1' after delay1 + 2177*delay_incr;
elsif nramp = '0' and StoredData = "100010000010" then SHout <= '1' after delay1 + 2178*delay_incr;
elsif nramp = '0' and StoredData = "100010000011" then SHout <= '1' after delay1 + 2179*delay_incr;
elsif nramp = '0' and StoredData = "100010000100" then SHout <= '1' after delay1 + 2180*delay_incr;
elsif nramp = '0' and StoredData = "100010000101" then SHout <= '1' after delay1 + 2181*delay_incr;
elsif nramp = '0' and StoredData = "100010000110" then SHout <= '1' after delay1 + 2182*delay_incr;
elsif nramp = '0' and StoredData = "100010000111" then SHout <= '1' after delay1 + 2183*delay_incr;
elsif nramp = '0' and StoredData = "100010001000" then SHout <= '1' after delay1 + 2184*delay_incr;
elsif nramp = '0' and StoredData = "100010001001" then SHout <= '1' after delay1 + 2185*delay_incr;
elsif nramp = '0' and StoredData = "100010001010" then SHout <= '1' after delay1 + 2186*delay_incr;
elsif nramp = '0' and StoredData = "100010001011" then SHout <= '1' after delay1 + 2187*delay_incr;
elsif nramp = '0' and StoredData = "100010001100" then SHout <= '1' after delay1 + 2188*delay_incr;
elsif nramp = '0' and StoredData = "100010001101" then SHout <= '1' after delay1 + 2189*delay_incr;
elsif nramp = '0' and StoredData = "100010001110" then SHout <= '1' after delay1 + 2190*delay_incr;
elsif nramp = '0' and StoredData = "100010001111" then SHout <= '1' after delay1 + 2191*delay_incr;
elsif nramp = '0' and StoredData = "100010010000" then SHout <= '1' after delay1 + 2192*delay_incr;
elsif nramp = '0' and StoredData = "100010010001" then SHout <= '1' after delay1 + 2193*delay_incr;
elsif nramp = '0' and StoredData = "100010010010" then SHout <= '1' after delay1 + 2194*delay_incr;
elsif nramp = '0' and StoredData = "100010010011" then SHout <= '1' after delay1 + 2195*delay_incr;
elsif nramp = '0' and StoredData = "100010010100" then SHout <= '1' after delay1 + 2196*delay_incr;
elsif nramp = '0' and StoredData = "100010010101" then SHout <= '1' after delay1 + 2197*delay_incr;
elsif nramp = '0' and StoredData = "100010010110" then SHout <= '1' after delay1 + 2198*delay_incr;
elsif nramp = '0' and StoredData = "100010010111" then SHout <= '1' after delay1 + 2199*delay_incr;
elsif nramp = '0' and StoredData = "100010011000" then SHout <= '1' after delay1 + 2200*delay_incr;
elsif nramp = '0' and StoredData = "100010011001" then SHout <= '1' after delay1 + 2201*delay_incr;
elsif nramp = '0' and StoredData = "100010011010" then SHout <= '1' after delay1 + 2202*delay_incr;
elsif nramp = '0' and StoredData = "100010011011" then SHout <= '1' after delay1 + 2203*delay_incr;
elsif nramp = '0' and StoredData = "100010011100" then SHout <= '1' after delay1 + 2204*delay_incr;
elsif nramp = '0' and StoredData = "100010011101" then SHout <= '1' after delay1 + 2205*delay_incr;
elsif nramp = '0' and StoredData = "100010011110" then SHout <= '1' after delay1 + 2206*delay_incr;
elsif nramp = '0' and StoredData = "100010011111" then SHout <= '1' after delay1 + 2207*delay_incr;
elsif nramp = '0' and StoredData = "100010100000" then SHout <= '1' after delay1 + 2208*delay_incr;
elsif nramp = '0' and StoredData = "100010100001" then SHout <= '1' after delay1 + 2209*delay_incr;
elsif nramp = '0' and StoredData = "100010100010" then SHout <= '1' after delay1 + 2210*delay_incr;
elsif nramp = '0' and StoredData = "100010100011" then SHout <= '1' after delay1 + 2211*delay_incr;
elsif nramp = '0' and StoredData = "100010100100" then SHout <= '1' after delay1 + 2212*delay_incr;
elsif nramp = '0' and StoredData = "100010100101" then SHout <= '1' after delay1 + 2213*delay_incr;
elsif nramp = '0' and StoredData = "100010100110" then SHout <= '1' after delay1 + 2214*delay_incr;
elsif nramp = '0' and StoredData = "100010100111" then SHout <= '1' after delay1 + 2215*delay_incr;
elsif nramp = '0' and StoredData = "100010101000" then SHout <= '1' after delay1 + 2216*delay_incr;
elsif nramp = '0' and StoredData = "100010101001" then SHout <= '1' after delay1 + 2217*delay_incr;
elsif nramp = '0' and StoredData = "100010101010" then SHout <= '1' after delay1 + 2218*delay_incr;
elsif nramp = '0' and StoredData = "100010101011" then SHout <= '1' after delay1 + 2219*delay_incr;
elsif nramp = '0' and StoredData = "100010101100" then SHout <= '1' after delay1 + 2220*delay_incr;
elsif nramp = '0' and StoredData = "100010101101" then SHout <= '1' after delay1 + 2221*delay_incr;
elsif nramp = '0' and StoredData = "100010101110" then SHout <= '1' after delay1 + 2222*delay_incr;
elsif nramp = '0' and StoredData = "100010101111" then SHout <= '1' after delay1 + 2223*delay_incr;
elsif nramp = '0' and StoredData = "100010110000" then SHout <= '1' after delay1 + 2224*delay_incr;
elsif nramp = '0' and StoredData = "100010110001" then SHout <= '1' after delay1 + 2225*delay_incr;
elsif nramp = '0' and StoredData = "100010110010" then SHout <= '1' after delay1 + 2226*delay_incr;
elsif nramp = '0' and StoredData = "100010110011" then SHout <= '1' after delay1 + 2227*delay_incr;
elsif nramp = '0' and StoredData = "100010110100" then SHout <= '1' after delay1 + 2228*delay_incr;
elsif nramp = '0' and StoredData = "100010110101" then SHout <= '1' after delay1 + 2229*delay_incr;
elsif nramp = '0' and StoredData = "100010110110" then SHout <= '1' after delay1 + 2230*delay_incr;
elsif nramp = '0' and StoredData = "100010110111" then SHout <= '1' after delay1 + 2231*delay_incr;
elsif nramp = '0' and StoredData = "100010111000" then SHout <= '1' after delay1 + 2232*delay_incr;
elsif nramp = '0' and StoredData = "100010111001" then SHout <= '1' after delay1 + 2233*delay_incr;
elsif nramp = '0' and StoredData = "100010111010" then SHout <= '1' after delay1 + 2234*delay_incr;
elsif nramp = '0' and StoredData = "100010111011" then SHout <= '1' after delay1 + 2235*delay_incr;
elsif nramp = '0' and StoredData = "100010111100" then SHout <= '1' after delay1 + 2236*delay_incr;
elsif nramp = '0' and StoredData = "100010111101" then SHout <= '1' after delay1 + 2237*delay_incr;
elsif nramp = '0' and StoredData = "100010111110" then SHout <= '1' after delay1 + 2238*delay_incr;
elsif nramp = '0' and StoredData = "100010111111" then SHout <= '1' after delay1 + 2239*delay_incr;
elsif nramp = '0' and StoredData = "100011000000" then SHout <= '1' after delay1 + 2240*delay_incr;
elsif nramp = '0' and StoredData = "100011000001" then SHout <= '1' after delay1 + 2241*delay_incr;
elsif nramp = '0' and StoredData = "100011000010" then SHout <= '1' after delay1 + 2242*delay_incr;
elsif nramp = '0' and StoredData = "100011000011" then SHout <= '1' after delay1 + 2243*delay_incr;
elsif nramp = '0' and StoredData = "100011000100" then SHout <= '1' after delay1 + 2244*delay_incr;
elsif nramp = '0' and StoredData = "100011000101" then SHout <= '1' after delay1 + 2245*delay_incr;
elsif nramp = '0' and StoredData = "100011000110" then SHout <= '1' after delay1 + 2246*delay_incr;
elsif nramp = '0' and StoredData = "100011000111" then SHout <= '1' after delay1 + 2247*delay_incr;
elsif nramp = '0' and StoredData = "100011001000" then SHout <= '1' after delay1 + 2248*delay_incr;
elsif nramp = '0' and StoredData = "100011001001" then SHout <= '1' after delay1 + 2249*delay_incr;
elsif nramp = '0' and StoredData = "100011001010" then SHout <= '1' after delay1 + 2250*delay_incr;
elsif nramp = '0' and StoredData = "100011001011" then SHout <= '1' after delay1 + 2251*delay_incr;
elsif nramp = '0' and StoredData = "100011001100" then SHout <= '1' after delay1 + 2252*delay_incr;
elsif nramp = '0' and StoredData = "100011001101" then SHout <= '1' after delay1 + 2253*delay_incr;
elsif nramp = '0' and StoredData = "100011001110" then SHout <= '1' after delay1 + 2254*delay_incr;
elsif nramp = '0' and StoredData = "100011001111" then SHout <= '1' after delay1 + 2255*delay_incr;
elsif nramp = '0' and StoredData = "100011010000" then SHout <= '1' after delay1 + 2256*delay_incr;
elsif nramp = '0' and StoredData = "100011010001" then SHout <= '1' after delay1 + 2257*delay_incr;
elsif nramp = '0' and StoredData = "100011010010" then SHout <= '1' after delay1 + 2258*delay_incr;
elsif nramp = '0' and StoredData = "100011010011" then SHout <= '1' after delay1 + 2259*delay_incr;
elsif nramp = '0' and StoredData = "100011010100" then SHout <= '1' after delay1 + 2260*delay_incr;
elsif nramp = '0' and StoredData = "100011010101" then SHout <= '1' after delay1 + 2261*delay_incr;
elsif nramp = '0' and StoredData = "100011010110" then SHout <= '1' after delay1 + 2262*delay_incr;
elsif nramp = '0' and StoredData = "100011010111" then SHout <= '1' after delay1 + 2263*delay_incr;
elsif nramp = '0' and StoredData = "100011011000" then SHout <= '1' after delay1 + 2264*delay_incr;
elsif nramp = '0' and StoredData = "100011011001" then SHout <= '1' after delay1 + 2265*delay_incr;
elsif nramp = '0' and StoredData = "100011011010" then SHout <= '1' after delay1 + 2266*delay_incr;
elsif nramp = '0' and StoredData = "100011011011" then SHout <= '1' after delay1 + 2267*delay_incr;
elsif nramp = '0' and StoredData = "100011011100" then SHout <= '1' after delay1 + 2268*delay_incr;
elsif nramp = '0' and StoredData = "100011011101" then SHout <= '1' after delay1 + 2269*delay_incr;
elsif nramp = '0' and StoredData = "100011011110" then SHout <= '1' after delay1 + 2270*delay_incr;
elsif nramp = '0' and StoredData = "100011011111" then SHout <= '1' after delay1 + 2271*delay_incr;
elsif nramp = '0' and StoredData = "100011100000" then SHout <= '1' after delay1 + 2272*delay_incr;
elsif nramp = '0' and StoredData = "100011100001" then SHout <= '1' after delay1 + 2273*delay_incr;
elsif nramp = '0' and StoredData = "100011100010" then SHout <= '1' after delay1 + 2274*delay_incr;
elsif nramp = '0' and StoredData = "100011100011" then SHout <= '1' after delay1 + 2275*delay_incr;
elsif nramp = '0' and StoredData = "100011100100" then SHout <= '1' after delay1 + 2276*delay_incr;
elsif nramp = '0' and StoredData = "100011100101" then SHout <= '1' after delay1 + 2277*delay_incr;
elsif nramp = '0' and StoredData = "100011100110" then SHout <= '1' after delay1 + 2278*delay_incr;
elsif nramp = '0' and StoredData = "100011100111" then SHout <= '1' after delay1 + 2279*delay_incr;
elsif nramp = '0' and StoredData = "100011101000" then SHout <= '1' after delay1 + 2280*delay_incr;
elsif nramp = '0' and StoredData = "100011101001" then SHout <= '1' after delay1 + 2281*delay_incr;
elsif nramp = '0' and StoredData = "100011101010" then SHout <= '1' after delay1 + 2282*delay_incr;
elsif nramp = '0' and StoredData = "100011101011" then SHout <= '1' after delay1 + 2283*delay_incr;
elsif nramp = '0' and StoredData = "100011101100" then SHout <= '1' after delay1 + 2284*delay_incr;
elsif nramp = '0' and StoredData = "100011101101" then SHout <= '1' after delay1 + 2285*delay_incr;
elsif nramp = '0' and StoredData = "100011101110" then SHout <= '1' after delay1 + 2286*delay_incr;
elsif nramp = '0' and StoredData = "100011101111" then SHout <= '1' after delay1 + 2287*delay_incr;
elsif nramp = '0' and StoredData = "100011110000" then SHout <= '1' after delay1 + 2288*delay_incr;
elsif nramp = '0' and StoredData = "100011110001" then SHout <= '1' after delay1 + 2289*delay_incr;
elsif nramp = '0' and StoredData = "100011110010" then SHout <= '1' after delay1 + 2290*delay_incr;
elsif nramp = '0' and StoredData = "100011110011" then SHout <= '1' after delay1 + 2291*delay_incr;
elsif nramp = '0' and StoredData = "100011110100" then SHout <= '1' after delay1 + 2292*delay_incr;
elsif nramp = '0' and StoredData = "100011110101" then SHout <= '1' after delay1 + 2293*delay_incr;
elsif nramp = '0' and StoredData = "100011110110" then SHout <= '1' after delay1 + 2294*delay_incr;
elsif nramp = '0' and StoredData = "100011110111" then SHout <= '1' after delay1 + 2295*delay_incr;
elsif nramp = '0' and StoredData = "100011111000" then SHout <= '1' after delay1 + 2296*delay_incr;
elsif nramp = '0' and StoredData = "100011111001" then SHout <= '1' after delay1 + 2297*delay_incr;
elsif nramp = '0' and StoredData = "100011111010" then SHout <= '1' after delay1 + 2298*delay_incr;
elsif nramp = '0' and StoredData = "100011111011" then SHout <= '1' after delay1 + 2299*delay_incr;
elsif nramp = '0' and StoredData = "100011111100" then SHout <= '1' after delay1 + 2300*delay_incr;
elsif nramp = '0' and StoredData = "100011111101" then SHout <= '1' after delay1 + 2301*delay_incr;
elsif nramp = '0' and StoredData = "100011111110" then SHout <= '1' after delay1 + 2302*delay_incr;
elsif nramp = '0' and StoredData = "100011111111" then SHout <= '1' after delay1 + 2303*delay_incr;
elsif nramp = '0' and StoredData = "100100000000" then SHout <= '1' after delay1 + 2304*delay_incr;
elsif nramp = '0' and StoredData = "100100000001" then SHout <= '1' after delay1 + 2305*delay_incr;
elsif nramp = '0' and StoredData = "100100000010" then SHout <= '1' after delay1 + 2306*delay_incr;
elsif nramp = '0' and StoredData = "100100000011" then SHout <= '1' after delay1 + 2307*delay_incr;
elsif nramp = '0' and StoredData = "100100000100" then SHout <= '1' after delay1 + 2308*delay_incr;
elsif nramp = '0' and StoredData = "100100000101" then SHout <= '1' after delay1 + 2309*delay_incr;
elsif nramp = '0' and StoredData = "100100000110" then SHout <= '1' after delay1 + 2310*delay_incr;
elsif nramp = '0' and StoredData = "100100000111" then SHout <= '1' after delay1 + 2311*delay_incr;
elsif nramp = '0' and StoredData = "100100001000" then SHout <= '1' after delay1 + 2312*delay_incr;
elsif nramp = '0' and StoredData = "100100001001" then SHout <= '1' after delay1 + 2313*delay_incr;
elsif nramp = '0' and StoredData = "100100001010" then SHout <= '1' after delay1 + 2314*delay_incr;
elsif nramp = '0' and StoredData = "100100001011" then SHout <= '1' after delay1 + 2315*delay_incr;
elsif nramp = '0' and StoredData = "100100001100" then SHout <= '1' after delay1 + 2316*delay_incr;
elsif nramp = '0' and StoredData = "100100001101" then SHout <= '1' after delay1 + 2317*delay_incr;
elsif nramp = '0' and StoredData = "100100001110" then SHout <= '1' after delay1 + 2318*delay_incr;
elsif nramp = '0' and StoredData = "100100001111" then SHout <= '1' after delay1 + 2319*delay_incr;
elsif nramp = '0' and StoredData = "100100010000" then SHout <= '1' after delay1 + 2320*delay_incr;
elsif nramp = '0' and StoredData = "100100010001" then SHout <= '1' after delay1 + 2321*delay_incr;
elsif nramp = '0' and StoredData = "100100010010" then SHout <= '1' after delay1 + 2322*delay_incr;
elsif nramp = '0' and StoredData = "100100010011" then SHout <= '1' after delay1 + 2323*delay_incr;
elsif nramp = '0' and StoredData = "100100010100" then SHout <= '1' after delay1 + 2324*delay_incr;
elsif nramp = '0' and StoredData = "100100010101" then SHout <= '1' after delay1 + 2325*delay_incr;
elsif nramp = '0' and StoredData = "100100010110" then SHout <= '1' after delay1 + 2326*delay_incr;
elsif nramp = '0' and StoredData = "100100010111" then SHout <= '1' after delay1 + 2327*delay_incr;
elsif nramp = '0' and StoredData = "100100011000" then SHout <= '1' after delay1 + 2328*delay_incr;
elsif nramp = '0' and StoredData = "100100011001" then SHout <= '1' after delay1 + 2329*delay_incr;
elsif nramp = '0' and StoredData = "100100011010" then SHout <= '1' after delay1 + 2330*delay_incr;
elsif nramp = '0' and StoredData = "100100011011" then SHout <= '1' after delay1 + 2331*delay_incr;
elsif nramp = '0' and StoredData = "100100011100" then SHout <= '1' after delay1 + 2332*delay_incr;
elsif nramp = '0' and StoredData = "100100011101" then SHout <= '1' after delay1 + 2333*delay_incr;
elsif nramp = '0' and StoredData = "100100011110" then SHout <= '1' after delay1 + 2334*delay_incr;
elsif nramp = '0' and StoredData = "100100011111" then SHout <= '1' after delay1 + 2335*delay_incr;
elsif nramp = '0' and StoredData = "100100100000" then SHout <= '1' after delay1 + 2336*delay_incr;
elsif nramp = '0' and StoredData = "100100100001" then SHout <= '1' after delay1 + 2337*delay_incr;
elsif nramp = '0' and StoredData = "100100100010" then SHout <= '1' after delay1 + 2338*delay_incr;
elsif nramp = '0' and StoredData = "100100100011" then SHout <= '1' after delay1 + 2339*delay_incr;
elsif nramp = '0' and StoredData = "100100100100" then SHout <= '1' after delay1 + 2340*delay_incr;
elsif nramp = '0' and StoredData = "100100100101" then SHout <= '1' after delay1 + 2341*delay_incr;
elsif nramp = '0' and StoredData = "100100100110" then SHout <= '1' after delay1 + 2342*delay_incr;
elsif nramp = '0' and StoredData = "100100100111" then SHout <= '1' after delay1 + 2343*delay_incr;
elsif nramp = '0' and StoredData = "100100101000" then SHout <= '1' after delay1 + 2344*delay_incr;
elsif nramp = '0' and StoredData = "100100101001" then SHout <= '1' after delay1 + 2345*delay_incr;
elsif nramp = '0' and StoredData = "100100101010" then SHout <= '1' after delay1 + 2346*delay_incr;
elsif nramp = '0' and StoredData = "100100101011" then SHout <= '1' after delay1 + 2347*delay_incr;
elsif nramp = '0' and StoredData = "100100101100" then SHout <= '1' after delay1 + 2348*delay_incr;
elsif nramp = '0' and StoredData = "100100101101" then SHout <= '1' after delay1 + 2349*delay_incr;
elsif nramp = '0' and StoredData = "100100101110" then SHout <= '1' after delay1 + 2350*delay_incr;
elsif nramp = '0' and StoredData = "100100101111" then SHout <= '1' after delay1 + 2351*delay_incr;
elsif nramp = '0' and StoredData = "100100110000" then SHout <= '1' after delay1 + 2352*delay_incr;
elsif nramp = '0' and StoredData = "100100110001" then SHout <= '1' after delay1 + 2353*delay_incr;
elsif nramp = '0' and StoredData = "100100110010" then SHout <= '1' after delay1 + 2354*delay_incr;
elsif nramp = '0' and StoredData = "100100110011" then SHout <= '1' after delay1 + 2355*delay_incr;
elsif nramp = '0' and StoredData = "100100110100" then SHout <= '1' after delay1 + 2356*delay_incr;
elsif nramp = '0' and StoredData = "100100110101" then SHout <= '1' after delay1 + 2357*delay_incr;
elsif nramp = '0' and StoredData = "100100110110" then SHout <= '1' after delay1 + 2358*delay_incr;
elsif nramp = '0' and StoredData = "100100110111" then SHout <= '1' after delay1 + 2359*delay_incr;
elsif nramp = '0' and StoredData = "100100111000" then SHout <= '1' after delay1 + 2360*delay_incr;
elsif nramp = '0' and StoredData = "100100111001" then SHout <= '1' after delay1 + 2361*delay_incr;
elsif nramp = '0' and StoredData = "100100111010" then SHout <= '1' after delay1 + 2362*delay_incr;
elsif nramp = '0' and StoredData = "100100111011" then SHout <= '1' after delay1 + 2363*delay_incr;
elsif nramp = '0' and StoredData = "100100111100" then SHout <= '1' after delay1 + 2364*delay_incr;
elsif nramp = '0' and StoredData = "100100111101" then SHout <= '1' after delay1 + 2365*delay_incr;
elsif nramp = '0' and StoredData = "100100111110" then SHout <= '1' after delay1 + 2366*delay_incr;
elsif nramp = '0' and StoredData = "100100111111" then SHout <= '1' after delay1 + 2367*delay_incr;
elsif nramp = '0' and StoredData = "100101000000" then SHout <= '1' after delay1 + 2368*delay_incr;
elsif nramp = '0' and StoredData = "100101000001" then SHout <= '1' after delay1 + 2369*delay_incr;
elsif nramp = '0' and StoredData = "100101000010" then SHout <= '1' after delay1 + 2370*delay_incr;
elsif nramp = '0' and StoredData = "100101000011" then SHout <= '1' after delay1 + 2371*delay_incr;
elsif nramp = '0' and StoredData = "100101000100" then SHout <= '1' after delay1 + 2372*delay_incr;
elsif nramp = '0' and StoredData = "100101000101" then SHout <= '1' after delay1 + 2373*delay_incr;
elsif nramp = '0' and StoredData = "100101000110" then SHout <= '1' after delay1 + 2374*delay_incr;
elsif nramp = '0' and StoredData = "100101000111" then SHout <= '1' after delay1 + 2375*delay_incr;
elsif nramp = '0' and StoredData = "100101001000" then SHout <= '1' after delay1 + 2376*delay_incr;
elsif nramp = '0' and StoredData = "100101001001" then SHout <= '1' after delay1 + 2377*delay_incr;
elsif nramp = '0' and StoredData = "100101001010" then SHout <= '1' after delay1 + 2378*delay_incr;
elsif nramp = '0' and StoredData = "100101001011" then SHout <= '1' after delay1 + 2379*delay_incr;
elsif nramp = '0' and StoredData = "100101001100" then SHout <= '1' after delay1 + 2380*delay_incr;
elsif nramp = '0' and StoredData = "100101001101" then SHout <= '1' after delay1 + 2381*delay_incr;
elsif nramp = '0' and StoredData = "100101001110" then SHout <= '1' after delay1 + 2382*delay_incr;
elsif nramp = '0' and StoredData = "100101001111" then SHout <= '1' after delay1 + 2383*delay_incr;
elsif nramp = '0' and StoredData = "100101010000" then SHout <= '1' after delay1 + 2384*delay_incr;
elsif nramp = '0' and StoredData = "100101010001" then SHout <= '1' after delay1 + 2385*delay_incr;
elsif nramp = '0' and StoredData = "100101010010" then SHout <= '1' after delay1 + 2386*delay_incr;
elsif nramp = '0' and StoredData = "100101010011" then SHout <= '1' after delay1 + 2387*delay_incr;
elsif nramp = '0' and StoredData = "100101010100" then SHout <= '1' after delay1 + 2388*delay_incr;
elsif nramp = '0' and StoredData = "100101010101" then SHout <= '1' after delay1 + 2389*delay_incr;
elsif nramp = '0' and StoredData = "100101010110" then SHout <= '1' after delay1 + 2390*delay_incr;
elsif nramp = '0' and StoredData = "100101010111" then SHout <= '1' after delay1 + 2391*delay_incr;
elsif nramp = '0' and StoredData = "100101011000" then SHout <= '1' after delay1 + 2392*delay_incr;
elsif nramp = '0' and StoredData = "100101011001" then SHout <= '1' after delay1 + 2393*delay_incr;
elsif nramp = '0' and StoredData = "100101011010" then SHout <= '1' after delay1 + 2394*delay_incr;
elsif nramp = '0' and StoredData = "100101011011" then SHout <= '1' after delay1 + 2395*delay_incr;
elsif nramp = '0' and StoredData = "100101011100" then SHout <= '1' after delay1 + 2396*delay_incr;
elsif nramp = '0' and StoredData = "100101011101" then SHout <= '1' after delay1 + 2397*delay_incr;
elsif nramp = '0' and StoredData = "100101011110" then SHout <= '1' after delay1 + 2398*delay_incr;
elsif nramp = '0' and StoredData = "100101011111" then SHout <= '1' after delay1 + 2399*delay_incr;
elsif nramp = '0' and StoredData = "100101100000" then SHout <= '1' after delay1 + 2400*delay_incr;
elsif nramp = '0' and StoredData = "100101100001" then SHout <= '1' after delay1 + 2401*delay_incr;
elsif nramp = '0' and StoredData = "100101100010" then SHout <= '1' after delay1 + 2402*delay_incr;
elsif nramp = '0' and StoredData = "100101100011" then SHout <= '1' after delay1 + 2403*delay_incr;
elsif nramp = '0' and StoredData = "100101100100" then SHout <= '1' after delay1 + 2404*delay_incr;
elsif nramp = '0' and StoredData = "100101100101" then SHout <= '1' after delay1 + 2405*delay_incr;
elsif nramp = '0' and StoredData = "100101100110" then SHout <= '1' after delay1 + 2406*delay_incr;
elsif nramp = '0' and StoredData = "100101100111" then SHout <= '1' after delay1 + 2407*delay_incr;
elsif nramp = '0' and StoredData = "100101101000" then SHout <= '1' after delay1 + 2408*delay_incr;
elsif nramp = '0' and StoredData = "100101101001" then SHout <= '1' after delay1 + 2409*delay_incr;
elsif nramp = '0' and StoredData = "100101101010" then SHout <= '1' after delay1 + 2410*delay_incr;
elsif nramp = '0' and StoredData = "100101101011" then SHout <= '1' after delay1 + 2411*delay_incr;
elsif nramp = '0' and StoredData = "100101101100" then SHout <= '1' after delay1 + 2412*delay_incr;
elsif nramp = '0' and StoredData = "100101101101" then SHout <= '1' after delay1 + 2413*delay_incr;
elsif nramp = '0' and StoredData = "100101101110" then SHout <= '1' after delay1 + 2414*delay_incr;
elsif nramp = '0' and StoredData = "100101101111" then SHout <= '1' after delay1 + 2415*delay_incr;
elsif nramp = '0' and StoredData = "100101110000" then SHout <= '1' after delay1 + 2416*delay_incr;
elsif nramp = '0' and StoredData = "100101110001" then SHout <= '1' after delay1 + 2417*delay_incr;
elsif nramp = '0' and StoredData = "100101110010" then SHout <= '1' after delay1 + 2418*delay_incr;
elsif nramp = '0' and StoredData = "100101110011" then SHout <= '1' after delay1 + 2419*delay_incr;
elsif nramp = '0' and StoredData = "100101110100" then SHout <= '1' after delay1 + 2420*delay_incr;
elsif nramp = '0' and StoredData = "100101110101" then SHout <= '1' after delay1 + 2421*delay_incr;
elsif nramp = '0' and StoredData = "100101110110" then SHout <= '1' after delay1 + 2422*delay_incr;
elsif nramp = '0' and StoredData = "100101110111" then SHout <= '1' after delay1 + 2423*delay_incr;
elsif nramp = '0' and StoredData = "100101111000" then SHout <= '1' after delay1 + 2424*delay_incr;
elsif nramp = '0' and StoredData = "100101111001" then SHout <= '1' after delay1 + 2425*delay_incr;
elsif nramp = '0' and StoredData = "100101111010" then SHout <= '1' after delay1 + 2426*delay_incr;
elsif nramp = '0' and StoredData = "100101111011" then SHout <= '1' after delay1 + 2427*delay_incr;
elsif nramp = '0' and StoredData = "100101111100" then SHout <= '1' after delay1 + 2428*delay_incr;
elsif nramp = '0' and StoredData = "100101111101" then SHout <= '1' after delay1 + 2429*delay_incr;
elsif nramp = '0' and StoredData = "100101111110" then SHout <= '1' after delay1 + 2430*delay_incr;
elsif nramp = '0' and StoredData = "100101111111" then SHout <= '1' after delay1 + 2431*delay_incr;
elsif nramp = '0' and StoredData = "100110000000" then SHout <= '1' after delay1 + 2432*delay_incr;
elsif nramp = '0' and StoredData = "100110000001" then SHout <= '1' after delay1 + 2433*delay_incr;
elsif nramp = '0' and StoredData = "100110000010" then SHout <= '1' after delay1 + 2434*delay_incr;
elsif nramp = '0' and StoredData = "100110000011" then SHout <= '1' after delay1 + 2435*delay_incr;
elsif nramp = '0' and StoredData = "100110000100" then SHout <= '1' after delay1 + 2436*delay_incr;
elsif nramp = '0' and StoredData = "100110000101" then SHout <= '1' after delay1 + 2437*delay_incr;
elsif nramp = '0' and StoredData = "100110000110" then SHout <= '1' after delay1 + 2438*delay_incr;
elsif nramp = '0' and StoredData = "100110000111" then SHout <= '1' after delay1 + 2439*delay_incr;
elsif nramp = '0' and StoredData = "100110001000" then SHout <= '1' after delay1 + 2440*delay_incr;
elsif nramp = '0' and StoredData = "100110001001" then SHout <= '1' after delay1 + 2441*delay_incr;
elsif nramp = '0' and StoredData = "100110001010" then SHout <= '1' after delay1 + 2442*delay_incr;
elsif nramp = '0' and StoredData = "100110001011" then SHout <= '1' after delay1 + 2443*delay_incr;
elsif nramp = '0' and StoredData = "100110001100" then SHout <= '1' after delay1 + 2444*delay_incr;
elsif nramp = '0' and StoredData = "100110001101" then SHout <= '1' after delay1 + 2445*delay_incr;
elsif nramp = '0' and StoredData = "100110001110" then SHout <= '1' after delay1 + 2446*delay_incr;
elsif nramp = '0' and StoredData = "100110001111" then SHout <= '1' after delay1 + 2447*delay_incr;
elsif nramp = '0' and StoredData = "100110010000" then SHout <= '1' after delay1 + 2448*delay_incr;
elsif nramp = '0' and StoredData = "100110010001" then SHout <= '1' after delay1 + 2449*delay_incr;
elsif nramp = '0' and StoredData = "100110010010" then SHout <= '1' after delay1 + 2450*delay_incr;
elsif nramp = '0' and StoredData = "100110010011" then SHout <= '1' after delay1 + 2451*delay_incr;
elsif nramp = '0' and StoredData = "100110010100" then SHout <= '1' after delay1 + 2452*delay_incr;
elsif nramp = '0' and StoredData = "100110010101" then SHout <= '1' after delay1 + 2453*delay_incr;
elsif nramp = '0' and StoredData = "100110010110" then SHout <= '1' after delay1 + 2454*delay_incr;
elsif nramp = '0' and StoredData = "100110010111" then SHout <= '1' after delay1 + 2455*delay_incr;
elsif nramp = '0' and StoredData = "100110011000" then SHout <= '1' after delay1 + 2456*delay_incr;
elsif nramp = '0' and StoredData = "100110011001" then SHout <= '1' after delay1 + 2457*delay_incr;
elsif nramp = '0' and StoredData = "100110011010" then SHout <= '1' after delay1 + 2458*delay_incr;
elsif nramp = '0' and StoredData = "100110011011" then SHout <= '1' after delay1 + 2459*delay_incr;
elsif nramp = '0' and StoredData = "100110011100" then SHout <= '1' after delay1 + 2460*delay_incr;
elsif nramp = '0' and StoredData = "100110011101" then SHout <= '1' after delay1 + 2461*delay_incr;
elsif nramp = '0' and StoredData = "100110011110" then SHout <= '1' after delay1 + 2462*delay_incr;
elsif nramp = '0' and StoredData = "100110011111" then SHout <= '1' after delay1 + 2463*delay_incr;
elsif nramp = '0' and StoredData = "100110100000" then SHout <= '1' after delay1 + 2464*delay_incr;
elsif nramp = '0' and StoredData = "100110100001" then SHout <= '1' after delay1 + 2465*delay_incr;
elsif nramp = '0' and StoredData = "100110100010" then SHout <= '1' after delay1 + 2466*delay_incr;
elsif nramp = '0' and StoredData = "100110100011" then SHout <= '1' after delay1 + 2467*delay_incr;
elsif nramp = '0' and StoredData = "100110100100" then SHout <= '1' after delay1 + 2468*delay_incr;
elsif nramp = '0' and StoredData = "100110100101" then SHout <= '1' after delay1 + 2469*delay_incr;
elsif nramp = '0' and StoredData = "100110100110" then SHout <= '1' after delay1 + 2470*delay_incr;
elsif nramp = '0' and StoredData = "100110100111" then SHout <= '1' after delay1 + 2471*delay_incr;
elsif nramp = '0' and StoredData = "100110101000" then SHout <= '1' after delay1 + 2472*delay_incr;
elsif nramp = '0' and StoredData = "100110101001" then SHout <= '1' after delay1 + 2473*delay_incr;
elsif nramp = '0' and StoredData = "100110101010" then SHout <= '1' after delay1 + 2474*delay_incr;
elsif nramp = '0' and StoredData = "100110101011" then SHout <= '1' after delay1 + 2475*delay_incr;
elsif nramp = '0' and StoredData = "100110101100" then SHout <= '1' after delay1 + 2476*delay_incr;
elsif nramp = '0' and StoredData = "100110101101" then SHout <= '1' after delay1 + 2477*delay_incr;
elsif nramp = '0' and StoredData = "100110101110" then SHout <= '1' after delay1 + 2478*delay_incr;
elsif nramp = '0' and StoredData = "100110101111" then SHout <= '1' after delay1 + 2479*delay_incr;
elsif nramp = '0' and StoredData = "100110110000" then SHout <= '1' after delay1 + 2480*delay_incr;
elsif nramp = '0' and StoredData = "100110110001" then SHout <= '1' after delay1 + 2481*delay_incr;
elsif nramp = '0' and StoredData = "100110110010" then SHout <= '1' after delay1 + 2482*delay_incr;
elsif nramp = '0' and StoredData = "100110110011" then SHout <= '1' after delay1 + 2483*delay_incr;
elsif nramp = '0' and StoredData = "100110110100" then SHout <= '1' after delay1 + 2484*delay_incr;
elsif nramp = '0' and StoredData = "100110110101" then SHout <= '1' after delay1 + 2485*delay_incr;
elsif nramp = '0' and StoredData = "100110110110" then SHout <= '1' after delay1 + 2486*delay_incr;
elsif nramp = '0' and StoredData = "100110110111" then SHout <= '1' after delay1 + 2487*delay_incr;
elsif nramp = '0' and StoredData = "100110111000" then SHout <= '1' after delay1 + 2488*delay_incr;
elsif nramp = '0' and StoredData = "100110111001" then SHout <= '1' after delay1 + 2489*delay_incr;
elsif nramp = '0' and StoredData = "100110111010" then SHout <= '1' after delay1 + 2490*delay_incr;
elsif nramp = '0' and StoredData = "100110111011" then SHout <= '1' after delay1 + 2491*delay_incr;
elsif nramp = '0' and StoredData = "100110111100" then SHout <= '1' after delay1 + 2492*delay_incr;
elsif nramp = '0' and StoredData = "100110111101" then SHout <= '1' after delay1 + 2493*delay_incr;
elsif nramp = '0' and StoredData = "100110111110" then SHout <= '1' after delay1 + 2494*delay_incr;
elsif nramp = '0' and StoredData = "100110111111" then SHout <= '1' after delay1 + 2495*delay_incr;
elsif nramp = '0' and StoredData = "100111000000" then SHout <= '1' after delay1 + 2496*delay_incr;
elsif nramp = '0' and StoredData = "100111000001" then SHout <= '1' after delay1 + 2497*delay_incr;
elsif nramp = '0' and StoredData = "100111000010" then SHout <= '1' after delay1 + 2498*delay_incr;
elsif nramp = '0' and StoredData = "100111000011" then SHout <= '1' after delay1 + 2499*delay_incr;
elsif nramp = '0' and StoredData = "100111000100" then SHout <= '1' after delay1 + 2500*delay_incr;
elsif nramp = '0' and StoredData = "100111000101" then SHout <= '1' after delay1 + 2501*delay_incr;
elsif nramp = '0' and StoredData = "100111000110" then SHout <= '1' after delay1 + 2502*delay_incr;
elsif nramp = '0' and StoredData = "100111000111" then SHout <= '1' after delay1 + 2503*delay_incr;
elsif nramp = '0' and StoredData = "100111001000" then SHout <= '1' after delay1 + 2504*delay_incr;
elsif nramp = '0' and StoredData = "100111001001" then SHout <= '1' after delay1 + 2505*delay_incr;
elsif nramp = '0' and StoredData = "100111001010" then SHout <= '1' after delay1 + 2506*delay_incr;
elsif nramp = '0' and StoredData = "100111001011" then SHout <= '1' after delay1 + 2507*delay_incr;
elsif nramp = '0' and StoredData = "100111001100" then SHout <= '1' after delay1 + 2508*delay_incr;
elsif nramp = '0' and StoredData = "100111001101" then SHout <= '1' after delay1 + 2509*delay_incr;
elsif nramp = '0' and StoredData = "100111001110" then SHout <= '1' after delay1 + 2510*delay_incr;
elsif nramp = '0' and StoredData = "100111001111" then SHout <= '1' after delay1 + 2511*delay_incr;
elsif nramp = '0' and StoredData = "100111010000" then SHout <= '1' after delay1 + 2512*delay_incr;
elsif nramp = '0' and StoredData = "100111010001" then SHout <= '1' after delay1 + 2513*delay_incr;
elsif nramp = '0' and StoredData = "100111010010" then SHout <= '1' after delay1 + 2514*delay_incr;
elsif nramp = '0' and StoredData = "100111010011" then SHout <= '1' after delay1 + 2515*delay_incr;
elsif nramp = '0' and StoredData = "100111010100" then SHout <= '1' after delay1 + 2516*delay_incr;
elsif nramp = '0' and StoredData = "100111010101" then SHout <= '1' after delay1 + 2517*delay_incr;
elsif nramp = '0' and StoredData = "100111010110" then SHout <= '1' after delay1 + 2518*delay_incr;
elsif nramp = '0' and StoredData = "100111010111" then SHout <= '1' after delay1 + 2519*delay_incr;
elsif nramp = '0' and StoredData = "100111011000" then SHout <= '1' after delay1 + 2520*delay_incr;
elsif nramp = '0' and StoredData = "100111011001" then SHout <= '1' after delay1 + 2521*delay_incr;
elsif nramp = '0' and StoredData = "100111011010" then SHout <= '1' after delay1 + 2522*delay_incr;
elsif nramp = '0' and StoredData = "100111011011" then SHout <= '1' after delay1 + 2523*delay_incr;
elsif nramp = '0' and StoredData = "100111011100" then SHout <= '1' after delay1 + 2524*delay_incr;
elsif nramp = '0' and StoredData = "100111011101" then SHout <= '1' after delay1 + 2525*delay_incr;
elsif nramp = '0' and StoredData = "100111011110" then SHout <= '1' after delay1 + 2526*delay_incr;
elsif nramp = '0' and StoredData = "100111011111" then SHout <= '1' after delay1 + 2527*delay_incr;
elsif nramp = '0' and StoredData = "100111100000" then SHout <= '1' after delay1 + 2528*delay_incr;
elsif nramp = '0' and StoredData = "100111100001" then SHout <= '1' after delay1 + 2529*delay_incr;
elsif nramp = '0' and StoredData = "100111100010" then SHout <= '1' after delay1 + 2530*delay_incr;
elsif nramp = '0' and StoredData = "100111100011" then SHout <= '1' after delay1 + 2531*delay_incr;
elsif nramp = '0' and StoredData = "100111100100" then SHout <= '1' after delay1 + 2532*delay_incr;
elsif nramp = '0' and StoredData = "100111100101" then SHout <= '1' after delay1 + 2533*delay_incr;
elsif nramp = '0' and StoredData = "100111100110" then SHout <= '1' after delay1 + 2534*delay_incr;
elsif nramp = '0' and StoredData = "100111100111" then SHout <= '1' after delay1 + 2535*delay_incr;
elsif nramp = '0' and StoredData = "100111101000" then SHout <= '1' after delay1 + 2536*delay_incr;
elsif nramp = '0' and StoredData = "100111101001" then SHout <= '1' after delay1 + 2537*delay_incr;
elsif nramp = '0' and StoredData = "100111101010" then SHout <= '1' after delay1 + 2538*delay_incr;
elsif nramp = '0' and StoredData = "100111101011" then SHout <= '1' after delay1 + 2539*delay_incr;
elsif nramp = '0' and StoredData = "100111101100" then SHout <= '1' after delay1 + 2540*delay_incr;
elsif nramp = '0' and StoredData = "100111101101" then SHout <= '1' after delay1 + 2541*delay_incr;
elsif nramp = '0' and StoredData = "100111101110" then SHout <= '1' after delay1 + 2542*delay_incr;
elsif nramp = '0' and StoredData = "100111101111" then SHout <= '1' after delay1 + 2543*delay_incr;
elsif nramp = '0' and StoredData = "100111110000" then SHout <= '1' after delay1 + 2544*delay_incr;
elsif nramp = '0' and StoredData = "100111110001" then SHout <= '1' after delay1 + 2545*delay_incr;
elsif nramp = '0' and StoredData = "100111110010" then SHout <= '1' after delay1 + 2546*delay_incr;
elsif nramp = '0' and StoredData = "100111110011" then SHout <= '1' after delay1 + 2547*delay_incr;
elsif nramp = '0' and StoredData = "100111110100" then SHout <= '1' after delay1 + 2548*delay_incr;
elsif nramp = '0' and StoredData = "100111110101" then SHout <= '1' after delay1 + 2549*delay_incr;
elsif nramp = '0' and StoredData = "100111110110" then SHout <= '1' after delay1 + 2550*delay_incr;
elsif nramp = '0' and StoredData = "100111110111" then SHout <= '1' after delay1 + 2551*delay_incr;
elsif nramp = '0' and StoredData = "100111111000" then SHout <= '1' after delay1 + 2552*delay_incr;
elsif nramp = '0' and StoredData = "100111111001" then SHout <= '1' after delay1 + 2553*delay_incr;
elsif nramp = '0' and StoredData = "100111111010" then SHout <= '1' after delay1 + 2554*delay_incr;
elsif nramp = '0' and StoredData = "100111111011" then SHout <= '1' after delay1 + 2555*delay_incr;
elsif nramp = '0' and StoredData = "100111111100" then SHout <= '1' after delay1 + 2556*delay_incr;
elsif nramp = '0' and StoredData = "100111111101" then SHout <= '1' after delay1 + 2557*delay_incr;
elsif nramp = '0' and StoredData = "100111111110" then SHout <= '1' after delay1 + 2558*delay_incr;
elsif nramp = '0' and StoredData = "100111111111" then SHout <= '1' after delay1 + 2559*delay_incr;
elsif nramp = '0' and StoredData = "101000000000" then SHout <= '1' after delay1 + 2560*delay_incr;
elsif nramp = '0' and StoredData = "101000000001" then SHout <= '1' after delay1 + 2561*delay_incr;
elsif nramp = '0' and StoredData = "101000000010" then SHout <= '1' after delay1 + 2562*delay_incr;
elsif nramp = '0' and StoredData = "101000000011" then SHout <= '1' after delay1 + 2563*delay_incr;
elsif nramp = '0' and StoredData = "101000000100" then SHout <= '1' after delay1 + 2564*delay_incr;
elsif nramp = '0' and StoredData = "101000000101" then SHout <= '1' after delay1 + 2565*delay_incr;
elsif nramp = '0' and StoredData = "101000000110" then SHout <= '1' after delay1 + 2566*delay_incr;
elsif nramp = '0' and StoredData = "101000000111" then SHout <= '1' after delay1 + 2567*delay_incr;
elsif nramp = '0' and StoredData = "101000001000" then SHout <= '1' after delay1 + 2568*delay_incr;
elsif nramp = '0' and StoredData = "101000001001" then SHout <= '1' after delay1 + 2569*delay_incr;
elsif nramp = '0' and StoredData = "101000001010" then SHout <= '1' after delay1 + 2570*delay_incr;
elsif nramp = '0' and StoredData = "101000001011" then SHout <= '1' after delay1 + 2571*delay_incr;
elsif nramp = '0' and StoredData = "101000001100" then SHout <= '1' after delay1 + 2572*delay_incr;
elsif nramp = '0' and StoredData = "101000001101" then SHout <= '1' after delay1 + 2573*delay_incr;
elsif nramp = '0' and StoredData = "101000001110" then SHout <= '1' after delay1 + 2574*delay_incr;
elsif nramp = '0' and StoredData = "101000001111" then SHout <= '1' after delay1 + 2575*delay_incr;
elsif nramp = '0' and StoredData = "101000010000" then SHout <= '1' after delay1 + 2576*delay_incr;
elsif nramp = '0' and StoredData = "101000010001" then SHout <= '1' after delay1 + 2577*delay_incr;
elsif nramp = '0' and StoredData = "101000010010" then SHout <= '1' after delay1 + 2578*delay_incr;
elsif nramp = '0' and StoredData = "101000010011" then SHout <= '1' after delay1 + 2579*delay_incr;
elsif nramp = '0' and StoredData = "101000010100" then SHout <= '1' after delay1 + 2580*delay_incr;
elsif nramp = '0' and StoredData = "101000010101" then SHout <= '1' after delay1 + 2581*delay_incr;
elsif nramp = '0' and StoredData = "101000010110" then SHout <= '1' after delay1 + 2582*delay_incr;
elsif nramp = '0' and StoredData = "101000010111" then SHout <= '1' after delay1 + 2583*delay_incr;
elsif nramp = '0' and StoredData = "101000011000" then SHout <= '1' after delay1 + 2584*delay_incr;
elsif nramp = '0' and StoredData = "101000011001" then SHout <= '1' after delay1 + 2585*delay_incr;
elsif nramp = '0' and StoredData = "101000011010" then SHout <= '1' after delay1 + 2586*delay_incr;
elsif nramp = '0' and StoredData = "101000011011" then SHout <= '1' after delay1 + 2587*delay_incr;
elsif nramp = '0' and StoredData = "101000011100" then SHout <= '1' after delay1 + 2588*delay_incr;
elsif nramp = '0' and StoredData = "101000011101" then SHout <= '1' after delay1 + 2589*delay_incr;
elsif nramp = '0' and StoredData = "101000011110" then SHout <= '1' after delay1 + 2590*delay_incr;
elsif nramp = '0' and StoredData = "101000011111" then SHout <= '1' after delay1 + 2591*delay_incr;
elsif nramp = '0' and StoredData = "101000100000" then SHout <= '1' after delay1 + 2592*delay_incr;
elsif nramp = '0' and StoredData = "101000100001" then SHout <= '1' after delay1 + 2593*delay_incr;
elsif nramp = '0' and StoredData = "101000100010" then SHout <= '1' after delay1 + 2594*delay_incr;
elsif nramp = '0' and StoredData = "101000100011" then SHout <= '1' after delay1 + 2595*delay_incr;
elsif nramp = '0' and StoredData = "101000100100" then SHout <= '1' after delay1 + 2596*delay_incr;
elsif nramp = '0' and StoredData = "101000100101" then SHout <= '1' after delay1 + 2597*delay_incr;
elsif nramp = '0' and StoredData = "101000100110" then SHout <= '1' after delay1 + 2598*delay_incr;
elsif nramp = '0' and StoredData = "101000100111" then SHout <= '1' after delay1 + 2599*delay_incr;
elsif nramp = '0' and StoredData = "101000101000" then SHout <= '1' after delay1 + 2600*delay_incr;
elsif nramp = '0' and StoredData = "101000101001" then SHout <= '1' after delay1 + 2601*delay_incr;
elsif nramp = '0' and StoredData = "101000101010" then SHout <= '1' after delay1 + 2602*delay_incr;
elsif nramp = '0' and StoredData = "101000101011" then SHout <= '1' after delay1 + 2603*delay_incr;
elsif nramp = '0' and StoredData = "101000101100" then SHout <= '1' after delay1 + 2604*delay_incr;
elsif nramp = '0' and StoredData = "101000101101" then SHout <= '1' after delay1 + 2605*delay_incr;
elsif nramp = '0' and StoredData = "101000101110" then SHout <= '1' after delay1 + 2606*delay_incr;
elsif nramp = '0' and StoredData = "101000101111" then SHout <= '1' after delay1 + 2607*delay_incr;
elsif nramp = '0' and StoredData = "101000110000" then SHout <= '1' after delay1 + 2608*delay_incr;
elsif nramp = '0' and StoredData = "101000110001" then SHout <= '1' after delay1 + 2609*delay_incr;
elsif nramp = '0' and StoredData = "101000110010" then SHout <= '1' after delay1 + 2610*delay_incr;
elsif nramp = '0' and StoredData = "101000110011" then SHout <= '1' after delay1 + 2611*delay_incr;
elsif nramp = '0' and StoredData = "101000110100" then SHout <= '1' after delay1 + 2612*delay_incr;
elsif nramp = '0' and StoredData = "101000110101" then SHout <= '1' after delay1 + 2613*delay_incr;
elsif nramp = '0' and StoredData = "101000110110" then SHout <= '1' after delay1 + 2614*delay_incr;
elsif nramp = '0' and StoredData = "101000110111" then SHout <= '1' after delay1 + 2615*delay_incr;
elsif nramp = '0' and StoredData = "101000111000" then SHout <= '1' after delay1 + 2616*delay_incr;
elsif nramp = '0' and StoredData = "101000111001" then SHout <= '1' after delay1 + 2617*delay_incr;
elsif nramp = '0' and StoredData = "101000111010" then SHout <= '1' after delay1 + 2618*delay_incr;
elsif nramp = '0' and StoredData = "101000111011" then SHout <= '1' after delay1 + 2619*delay_incr;
elsif nramp = '0' and StoredData = "101000111100" then SHout <= '1' after delay1 + 2620*delay_incr;
elsif nramp = '0' and StoredData = "101000111101" then SHout <= '1' after delay1 + 2621*delay_incr;
elsif nramp = '0' and StoredData = "101000111110" then SHout <= '1' after delay1 + 2622*delay_incr;
elsif nramp = '0' and StoredData = "101000111111" then SHout <= '1' after delay1 + 2623*delay_incr;
elsif nramp = '0' and StoredData = "101001000000" then SHout <= '1' after delay1 + 2624*delay_incr;
elsif nramp = '0' and StoredData = "101001000001" then SHout <= '1' after delay1 + 2625*delay_incr;
elsif nramp = '0' and StoredData = "101001000010" then SHout <= '1' after delay1 + 2626*delay_incr;
elsif nramp = '0' and StoredData = "101001000011" then SHout <= '1' after delay1 + 2627*delay_incr;
elsif nramp = '0' and StoredData = "101001000100" then SHout <= '1' after delay1 + 2628*delay_incr;
elsif nramp = '0' and StoredData = "101001000101" then SHout <= '1' after delay1 + 2629*delay_incr;
elsif nramp = '0' and StoredData = "101001000110" then SHout <= '1' after delay1 + 2630*delay_incr;
elsif nramp = '0' and StoredData = "101001000111" then SHout <= '1' after delay1 + 2631*delay_incr;
elsif nramp = '0' and StoredData = "101001001000" then SHout <= '1' after delay1 + 2632*delay_incr;
elsif nramp = '0' and StoredData = "101001001001" then SHout <= '1' after delay1 + 2633*delay_incr;
elsif nramp = '0' and StoredData = "101001001010" then SHout <= '1' after delay1 + 2634*delay_incr;
elsif nramp = '0' and StoredData = "101001001011" then SHout <= '1' after delay1 + 2635*delay_incr;
elsif nramp = '0' and StoredData = "101001001100" then SHout <= '1' after delay1 + 2636*delay_incr;
elsif nramp = '0' and StoredData = "101001001101" then SHout <= '1' after delay1 + 2637*delay_incr;
elsif nramp = '0' and StoredData = "101001001110" then SHout <= '1' after delay1 + 2638*delay_incr;
elsif nramp = '0' and StoredData = "101001001111" then SHout <= '1' after delay1 + 2639*delay_incr;
elsif nramp = '0' and StoredData = "101001010000" then SHout <= '1' after delay1 + 2640*delay_incr;
elsif nramp = '0' and StoredData = "101001010001" then SHout <= '1' after delay1 + 2641*delay_incr;
elsif nramp = '0' and StoredData = "101001010010" then SHout <= '1' after delay1 + 2642*delay_incr;
elsif nramp = '0' and StoredData = "101001010011" then SHout <= '1' after delay1 + 2643*delay_incr;
elsif nramp = '0' and StoredData = "101001010100" then SHout <= '1' after delay1 + 2644*delay_incr;
elsif nramp = '0' and StoredData = "101001010101" then SHout <= '1' after delay1 + 2645*delay_incr;
elsif nramp = '0' and StoredData = "101001010110" then SHout <= '1' after delay1 + 2646*delay_incr;
elsif nramp = '0' and StoredData = "101001010111" then SHout <= '1' after delay1 + 2647*delay_incr;
elsif nramp = '0' and StoredData = "101001011000" then SHout <= '1' after delay1 + 2648*delay_incr;
elsif nramp = '0' and StoredData = "101001011001" then SHout <= '1' after delay1 + 2649*delay_incr;
elsif nramp = '0' and StoredData = "101001011010" then SHout <= '1' after delay1 + 2650*delay_incr;
elsif nramp = '0' and StoredData = "101001011011" then SHout <= '1' after delay1 + 2651*delay_incr;
elsif nramp = '0' and StoredData = "101001011100" then SHout <= '1' after delay1 + 2652*delay_incr;
elsif nramp = '0' and StoredData = "101001011101" then SHout <= '1' after delay1 + 2653*delay_incr;
elsif nramp = '0' and StoredData = "101001011110" then SHout <= '1' after delay1 + 2654*delay_incr;
elsif nramp = '0' and StoredData = "101001011111" then SHout <= '1' after delay1 + 2655*delay_incr;
elsif nramp = '0' and StoredData = "101001100000" then SHout <= '1' after delay1 + 2656*delay_incr;
elsif nramp = '0' and StoredData = "101001100001" then SHout <= '1' after delay1 + 2657*delay_incr;
elsif nramp = '0' and StoredData = "101001100010" then SHout <= '1' after delay1 + 2658*delay_incr;
elsif nramp = '0' and StoredData = "101001100011" then SHout <= '1' after delay1 + 2659*delay_incr;
elsif nramp = '0' and StoredData = "101001100100" then SHout <= '1' after delay1 + 2660*delay_incr;
elsif nramp = '0' and StoredData = "101001100101" then SHout <= '1' after delay1 + 2661*delay_incr;
elsif nramp = '0' and StoredData = "101001100110" then SHout <= '1' after delay1 + 2662*delay_incr;
elsif nramp = '0' and StoredData = "101001100111" then SHout <= '1' after delay1 + 2663*delay_incr;
elsif nramp = '0' and StoredData = "101001101000" then SHout <= '1' after delay1 + 2664*delay_incr;
elsif nramp = '0' and StoredData = "101001101001" then SHout <= '1' after delay1 + 2665*delay_incr;
elsif nramp = '0' and StoredData = "101001101010" then SHout <= '1' after delay1 + 2666*delay_incr;
elsif nramp = '0' and StoredData = "101001101011" then SHout <= '1' after delay1 + 2667*delay_incr;
elsif nramp = '0' and StoredData = "101001101100" then SHout <= '1' after delay1 + 2668*delay_incr;
elsif nramp = '0' and StoredData = "101001101101" then SHout <= '1' after delay1 + 2669*delay_incr;
elsif nramp = '0' and StoredData = "101001101110" then SHout <= '1' after delay1 + 2670*delay_incr;
elsif nramp = '0' and StoredData = "101001101111" then SHout <= '1' after delay1 + 2671*delay_incr;
elsif nramp = '0' and StoredData = "101001110000" then SHout <= '1' after delay1 + 2672*delay_incr;
elsif nramp = '0' and StoredData = "101001110001" then SHout <= '1' after delay1 + 2673*delay_incr;
elsif nramp = '0' and StoredData = "101001110010" then SHout <= '1' after delay1 + 2674*delay_incr;
elsif nramp = '0' and StoredData = "101001110011" then SHout <= '1' after delay1 + 2675*delay_incr;
elsif nramp = '0' and StoredData = "101001110100" then SHout <= '1' after delay1 + 2676*delay_incr;
elsif nramp = '0' and StoredData = "101001110101" then SHout <= '1' after delay1 + 2677*delay_incr;
elsif nramp = '0' and StoredData = "101001110110" then SHout <= '1' after delay1 + 2678*delay_incr;
elsif nramp = '0' and StoredData = "101001110111" then SHout <= '1' after delay1 + 2679*delay_incr;
elsif nramp = '0' and StoredData = "101001111000" then SHout <= '1' after delay1 + 2680*delay_incr;
elsif nramp = '0' and StoredData = "101001111001" then SHout <= '1' after delay1 + 2681*delay_incr;
elsif nramp = '0' and StoredData = "101001111010" then SHout <= '1' after delay1 + 2682*delay_incr;
elsif nramp = '0' and StoredData = "101001111011" then SHout <= '1' after delay1 + 2683*delay_incr;
elsif nramp = '0' and StoredData = "101001111100" then SHout <= '1' after delay1 + 2684*delay_incr;
elsif nramp = '0' and StoredData = "101001111101" then SHout <= '1' after delay1 + 2685*delay_incr;
elsif nramp = '0' and StoredData = "101001111110" then SHout <= '1' after delay1 + 2686*delay_incr;
elsif nramp = '0' and StoredData = "101001111111" then SHout <= '1' after delay1 + 2687*delay_incr;
elsif nramp = '0' and StoredData = "101010000000" then SHout <= '1' after delay1 + 2688*delay_incr;
elsif nramp = '0' and StoredData = "101010000001" then SHout <= '1' after delay1 + 2689*delay_incr;
elsif nramp = '0' and StoredData = "101010000010" then SHout <= '1' after delay1 + 2690*delay_incr;
elsif nramp = '0' and StoredData = "101010000011" then SHout <= '1' after delay1 + 2691*delay_incr;
elsif nramp = '0' and StoredData = "101010000100" then SHout <= '1' after delay1 + 2692*delay_incr;
elsif nramp = '0' and StoredData = "101010000101" then SHout <= '1' after delay1 + 2693*delay_incr;
elsif nramp = '0' and StoredData = "101010000110" then SHout <= '1' after delay1 + 2694*delay_incr;
elsif nramp = '0' and StoredData = "101010000111" then SHout <= '1' after delay1 + 2695*delay_incr;
elsif nramp = '0' and StoredData = "101010001000" then SHout <= '1' after delay1 + 2696*delay_incr;
elsif nramp = '0' and StoredData = "101010001001" then SHout <= '1' after delay1 + 2697*delay_incr;
elsif nramp = '0' and StoredData = "101010001010" then SHout <= '1' after delay1 + 2698*delay_incr;
elsif nramp = '0' and StoredData = "101010001011" then SHout <= '1' after delay1 + 2699*delay_incr;
elsif nramp = '0' and StoredData = "101010001100" then SHout <= '1' after delay1 + 2700*delay_incr;
elsif nramp = '0' and StoredData = "101010001101" then SHout <= '1' after delay1 + 2701*delay_incr;
elsif nramp = '0' and StoredData = "101010001110" then SHout <= '1' after delay1 + 2702*delay_incr;
elsif nramp = '0' and StoredData = "101010001111" then SHout <= '1' after delay1 + 2703*delay_incr;
elsif nramp = '0' and StoredData = "101010010000" then SHout <= '1' after delay1 + 2704*delay_incr;
elsif nramp = '0' and StoredData = "101010010001" then SHout <= '1' after delay1 + 2705*delay_incr;
elsif nramp = '0' and StoredData = "101010010010" then SHout <= '1' after delay1 + 2706*delay_incr;
elsif nramp = '0' and StoredData = "101010010011" then SHout <= '1' after delay1 + 2707*delay_incr;
elsif nramp = '0' and StoredData = "101010010100" then SHout <= '1' after delay1 + 2708*delay_incr;
elsif nramp = '0' and StoredData = "101010010101" then SHout <= '1' after delay1 + 2709*delay_incr;
elsif nramp = '0' and StoredData = "101010010110" then SHout <= '1' after delay1 + 2710*delay_incr;
elsif nramp = '0' and StoredData = "101010010111" then SHout <= '1' after delay1 + 2711*delay_incr;
elsif nramp = '0' and StoredData = "101010011000" then SHout <= '1' after delay1 + 2712*delay_incr;
elsif nramp = '0' and StoredData = "101010011001" then SHout <= '1' after delay1 + 2713*delay_incr;
elsif nramp = '0' and StoredData = "101010011010" then SHout <= '1' after delay1 + 2714*delay_incr;
elsif nramp = '0' and StoredData = "101010011011" then SHout <= '1' after delay1 + 2715*delay_incr;
elsif nramp = '0' and StoredData = "101010011100" then SHout <= '1' after delay1 + 2716*delay_incr;
elsif nramp = '0' and StoredData = "101010011101" then SHout <= '1' after delay1 + 2717*delay_incr;
elsif nramp = '0' and StoredData = "101010011110" then SHout <= '1' after delay1 + 2718*delay_incr;
elsif nramp = '0' and StoredData = "101010011111" then SHout <= '1' after delay1 + 2719*delay_incr;
elsif nramp = '0' and StoredData = "101010100000" then SHout <= '1' after delay1 + 2720*delay_incr;
elsif nramp = '0' and StoredData = "101010100001" then SHout <= '1' after delay1 + 2721*delay_incr;
elsif nramp = '0' and StoredData = "101010100010" then SHout <= '1' after delay1 + 2722*delay_incr;
elsif nramp = '0' and StoredData = "101010100011" then SHout <= '1' after delay1 + 2723*delay_incr;
elsif nramp = '0' and StoredData = "101010100100" then SHout <= '1' after delay1 + 2724*delay_incr;
elsif nramp = '0' and StoredData = "101010100101" then SHout <= '1' after delay1 + 2725*delay_incr;
elsif nramp = '0' and StoredData = "101010100110" then SHout <= '1' after delay1 + 2726*delay_incr;
elsif nramp = '0' and StoredData = "101010100111" then SHout <= '1' after delay1 + 2727*delay_incr;
elsif nramp = '0' and StoredData = "101010101000" then SHout <= '1' after delay1 + 2728*delay_incr;
elsif nramp = '0' and StoredData = "101010101001" then SHout <= '1' after delay1 + 2729*delay_incr;
elsif nramp = '0' and StoredData = "101010101010" then SHout <= '1' after delay1 + 2730*delay_incr;
elsif nramp = '0' and StoredData = "101010101011" then SHout <= '1' after delay1 + 2731*delay_incr;
elsif nramp = '0' and StoredData = "101010101100" then SHout <= '1' after delay1 + 2732*delay_incr;
elsif nramp = '0' and StoredData = "101010101101" then SHout <= '1' after delay1 + 2733*delay_incr;
elsif nramp = '0' and StoredData = "101010101110" then SHout <= '1' after delay1 + 2734*delay_incr;
elsif nramp = '0' and StoredData = "101010101111" then SHout <= '1' after delay1 + 2735*delay_incr;
elsif nramp = '0' and StoredData = "101010110000" then SHout <= '1' after delay1 + 2736*delay_incr;
elsif nramp = '0' and StoredData = "101010110001" then SHout <= '1' after delay1 + 2737*delay_incr;
elsif nramp = '0' and StoredData = "101010110010" then SHout <= '1' after delay1 + 2738*delay_incr;
elsif nramp = '0' and StoredData = "101010110011" then SHout <= '1' after delay1 + 2739*delay_incr;
elsif nramp = '0' and StoredData = "101010110100" then SHout <= '1' after delay1 + 2740*delay_incr;
elsif nramp = '0' and StoredData = "101010110101" then SHout <= '1' after delay1 + 2741*delay_incr;
elsif nramp = '0' and StoredData = "101010110110" then SHout <= '1' after delay1 + 2742*delay_incr;
elsif nramp = '0' and StoredData = "101010110111" then SHout <= '1' after delay1 + 2743*delay_incr;
elsif nramp = '0' and StoredData = "101010111000" then SHout <= '1' after delay1 + 2744*delay_incr;
elsif nramp = '0' and StoredData = "101010111001" then SHout <= '1' after delay1 + 2745*delay_incr;
elsif nramp = '0' and StoredData = "101010111010" then SHout <= '1' after delay1 + 2746*delay_incr;
elsif nramp = '0' and StoredData = "101010111011" then SHout <= '1' after delay1 + 2747*delay_incr;
elsif nramp = '0' and StoredData = "101010111100" then SHout <= '1' after delay1 + 2748*delay_incr;
elsif nramp = '0' and StoredData = "101010111101" then SHout <= '1' after delay1 + 2749*delay_incr;
elsif nramp = '0' and StoredData = "101010111110" then SHout <= '1' after delay1 + 2750*delay_incr;
elsif nramp = '0' and StoredData = "101010111111" then SHout <= '1' after delay1 + 2751*delay_incr;
elsif nramp = '0' and StoredData = "101011000000" then SHout <= '1' after delay1 + 2752*delay_incr;
elsif nramp = '0' and StoredData = "101011000001" then SHout <= '1' after delay1 + 2753*delay_incr;
elsif nramp = '0' and StoredData = "101011000010" then SHout <= '1' after delay1 + 2754*delay_incr;
elsif nramp = '0' and StoredData = "101011000011" then SHout <= '1' after delay1 + 2755*delay_incr;
elsif nramp = '0' and StoredData = "101011000100" then SHout <= '1' after delay1 + 2756*delay_incr;
elsif nramp = '0' and StoredData = "101011000101" then SHout <= '1' after delay1 + 2757*delay_incr;
elsif nramp = '0' and StoredData = "101011000110" then SHout <= '1' after delay1 + 2758*delay_incr;
elsif nramp = '0' and StoredData = "101011000111" then SHout <= '1' after delay1 + 2759*delay_incr;
elsif nramp = '0' and StoredData = "101011001000" then SHout <= '1' after delay1 + 2760*delay_incr;
elsif nramp = '0' and StoredData = "101011001001" then SHout <= '1' after delay1 + 2761*delay_incr;
elsif nramp = '0' and StoredData = "101011001010" then SHout <= '1' after delay1 + 2762*delay_incr;
elsif nramp = '0' and StoredData = "101011001011" then SHout <= '1' after delay1 + 2763*delay_incr;
elsif nramp = '0' and StoredData = "101011001100" then SHout <= '1' after delay1 + 2764*delay_incr;
elsif nramp = '0' and StoredData = "101011001101" then SHout <= '1' after delay1 + 2765*delay_incr;
elsif nramp = '0' and StoredData = "101011001110" then SHout <= '1' after delay1 + 2766*delay_incr;
elsif nramp = '0' and StoredData = "101011001111" then SHout <= '1' after delay1 + 2767*delay_incr;
elsif nramp = '0' and StoredData = "101011010000" then SHout <= '1' after delay1 + 2768*delay_incr;
elsif nramp = '0' and StoredData = "101011010001" then SHout <= '1' after delay1 + 2769*delay_incr;
elsif nramp = '0' and StoredData = "101011010010" then SHout <= '1' after delay1 + 2770*delay_incr;
elsif nramp = '0' and StoredData = "101011010011" then SHout <= '1' after delay1 + 2771*delay_incr;
elsif nramp = '0' and StoredData = "101011010100" then SHout <= '1' after delay1 + 2772*delay_incr;
elsif nramp = '0' and StoredData = "101011010101" then SHout <= '1' after delay1 + 2773*delay_incr;
elsif nramp = '0' and StoredData = "101011010110" then SHout <= '1' after delay1 + 2774*delay_incr;
elsif nramp = '0' and StoredData = "101011010111" then SHout <= '1' after delay1 + 2775*delay_incr;
elsif nramp = '0' and StoredData = "101011011000" then SHout <= '1' after delay1 + 2776*delay_incr;
elsif nramp = '0' and StoredData = "101011011001" then SHout <= '1' after delay1 + 2777*delay_incr;
elsif nramp = '0' and StoredData = "101011011010" then SHout <= '1' after delay1 + 2778*delay_incr;
elsif nramp = '0' and StoredData = "101011011011" then SHout <= '1' after delay1 + 2779*delay_incr;
elsif nramp = '0' and StoredData = "101011011100" then SHout <= '1' after delay1 + 2780*delay_incr;
elsif nramp = '0' and StoredData = "101011011101" then SHout <= '1' after delay1 + 2781*delay_incr;
elsif nramp = '0' and StoredData = "101011011110" then SHout <= '1' after delay1 + 2782*delay_incr;
elsif nramp = '0' and StoredData = "101011011111" then SHout <= '1' after delay1 + 2783*delay_incr;
elsif nramp = '0' and StoredData = "101011100000" then SHout <= '1' after delay1 + 2784*delay_incr;
elsif nramp = '0' and StoredData = "101011100001" then SHout <= '1' after delay1 + 2785*delay_incr;
elsif nramp = '0' and StoredData = "101011100010" then SHout <= '1' after delay1 + 2786*delay_incr;
elsif nramp = '0' and StoredData = "101011100011" then SHout <= '1' after delay1 + 2787*delay_incr;
elsif nramp = '0' and StoredData = "101011100100" then SHout <= '1' after delay1 + 2788*delay_incr;
elsif nramp = '0' and StoredData = "101011100101" then SHout <= '1' after delay1 + 2789*delay_incr;
elsif nramp = '0' and StoredData = "101011100110" then SHout <= '1' after delay1 + 2790*delay_incr;
elsif nramp = '0' and StoredData = "101011100111" then SHout <= '1' after delay1 + 2791*delay_incr;
elsif nramp = '0' and StoredData = "101011101000" then SHout <= '1' after delay1 + 2792*delay_incr;
elsif nramp = '0' and StoredData = "101011101001" then SHout <= '1' after delay1 + 2793*delay_incr;
elsif nramp = '0' and StoredData = "101011101010" then SHout <= '1' after delay1 + 2794*delay_incr;
elsif nramp = '0' and StoredData = "101011101011" then SHout <= '1' after delay1 + 2795*delay_incr;
elsif nramp = '0' and StoredData = "101011101100" then SHout <= '1' after delay1 + 2796*delay_incr;
elsif nramp = '0' and StoredData = "101011101101" then SHout <= '1' after delay1 + 2797*delay_incr;
elsif nramp = '0' and StoredData = "101011101110" then SHout <= '1' after delay1 + 2798*delay_incr;
elsif nramp = '0' and StoredData = "101011101111" then SHout <= '1' after delay1 + 2799*delay_incr;
elsif nramp = '0' and StoredData = "101011110000" then SHout <= '1' after delay1 + 2800*delay_incr;
elsif nramp = '0' and StoredData = "101011110001" then SHout <= '1' after delay1 + 2801*delay_incr;
elsif nramp = '0' and StoredData = "101011110010" then SHout <= '1' after delay1 + 2802*delay_incr;
elsif nramp = '0' and StoredData = "101011110011" then SHout <= '1' after delay1 + 2803*delay_incr;
elsif nramp = '0' and StoredData = "101011110100" then SHout <= '1' after delay1 + 2804*delay_incr;
elsif nramp = '0' and StoredData = "101011110101" then SHout <= '1' after delay1 + 2805*delay_incr;
elsif nramp = '0' and StoredData = "101011110110" then SHout <= '1' after delay1 + 2806*delay_incr;
elsif nramp = '0' and StoredData = "101011110111" then SHout <= '1' after delay1 + 2807*delay_incr;
elsif nramp = '0' and StoredData = "101011111000" then SHout <= '1' after delay1 + 2808*delay_incr;
elsif nramp = '0' and StoredData = "101011111001" then SHout <= '1' after delay1 + 2809*delay_incr;
elsif nramp = '0' and StoredData = "101011111010" then SHout <= '1' after delay1 + 2810*delay_incr;
elsif nramp = '0' and StoredData = "101011111011" then SHout <= '1' after delay1 + 2811*delay_incr;
elsif nramp = '0' and StoredData = "101011111100" then SHout <= '1' after delay1 + 2812*delay_incr;
elsif nramp = '0' and StoredData = "101011111101" then SHout <= '1' after delay1 + 2813*delay_incr;
elsif nramp = '0' and StoredData = "101011111110" then SHout <= '1' after delay1 + 2814*delay_incr;
elsif nramp = '0' and StoredData = "101011111111" then SHout <= '1' after delay1 + 2815*delay_incr;
elsif nramp = '0' and StoredData = "101100000000" then SHout <= '1' after delay1 + 2816*delay_incr;
elsif nramp = '0' and StoredData = "101100000001" then SHout <= '1' after delay1 + 2817*delay_incr;
elsif nramp = '0' and StoredData = "101100000010" then SHout <= '1' after delay1 + 2818*delay_incr;
elsif nramp = '0' and StoredData = "101100000011" then SHout <= '1' after delay1 + 2819*delay_incr;
elsif nramp = '0' and StoredData = "101100000100" then SHout <= '1' after delay1 + 2820*delay_incr;
elsif nramp = '0' and StoredData = "101100000101" then SHout <= '1' after delay1 + 2821*delay_incr;
elsif nramp = '0' and StoredData = "101100000110" then SHout <= '1' after delay1 + 2822*delay_incr;
elsif nramp = '0' and StoredData = "101100000111" then SHout <= '1' after delay1 + 2823*delay_incr;
elsif nramp = '0' and StoredData = "101100001000" then SHout <= '1' after delay1 + 2824*delay_incr;
elsif nramp = '0' and StoredData = "101100001001" then SHout <= '1' after delay1 + 2825*delay_incr;
elsif nramp = '0' and StoredData = "101100001010" then SHout <= '1' after delay1 + 2826*delay_incr;
elsif nramp = '0' and StoredData = "101100001011" then SHout <= '1' after delay1 + 2827*delay_incr;
elsif nramp = '0' and StoredData = "101100001100" then SHout <= '1' after delay1 + 2828*delay_incr;
elsif nramp = '0' and StoredData = "101100001101" then SHout <= '1' after delay1 + 2829*delay_incr;
elsif nramp = '0' and StoredData = "101100001110" then SHout <= '1' after delay1 + 2830*delay_incr;
elsif nramp = '0' and StoredData = "101100001111" then SHout <= '1' after delay1 + 2831*delay_incr;
elsif nramp = '0' and StoredData = "101100010000" then SHout <= '1' after delay1 + 2832*delay_incr;
elsif nramp = '0' and StoredData = "101100010001" then SHout <= '1' after delay1 + 2833*delay_incr;
elsif nramp = '0' and StoredData = "101100010010" then SHout <= '1' after delay1 + 2834*delay_incr;
elsif nramp = '0' and StoredData = "101100010011" then SHout <= '1' after delay1 + 2835*delay_incr;
elsif nramp = '0' and StoredData = "101100010100" then SHout <= '1' after delay1 + 2836*delay_incr;
elsif nramp = '0' and StoredData = "101100010101" then SHout <= '1' after delay1 + 2837*delay_incr;
elsif nramp = '0' and StoredData = "101100010110" then SHout <= '1' after delay1 + 2838*delay_incr;
elsif nramp = '0' and StoredData = "101100010111" then SHout <= '1' after delay1 + 2839*delay_incr;
elsif nramp = '0' and StoredData = "101100011000" then SHout <= '1' after delay1 + 2840*delay_incr;
elsif nramp = '0' and StoredData = "101100011001" then SHout <= '1' after delay1 + 2841*delay_incr;
elsif nramp = '0' and StoredData = "101100011010" then SHout <= '1' after delay1 + 2842*delay_incr;
elsif nramp = '0' and StoredData = "101100011011" then SHout <= '1' after delay1 + 2843*delay_incr;
elsif nramp = '0' and StoredData = "101100011100" then SHout <= '1' after delay1 + 2844*delay_incr;
elsif nramp = '0' and StoredData = "101100011101" then SHout <= '1' after delay1 + 2845*delay_incr;
elsif nramp = '0' and StoredData = "101100011110" then SHout <= '1' after delay1 + 2846*delay_incr;
elsif nramp = '0' and StoredData = "101100011111" then SHout <= '1' after delay1 + 2847*delay_incr;
elsif nramp = '0' and StoredData = "101100100000" then SHout <= '1' after delay1 + 2848*delay_incr;
elsif nramp = '0' and StoredData = "101100100001" then SHout <= '1' after delay1 + 2849*delay_incr;
elsif nramp = '0' and StoredData = "101100100010" then SHout <= '1' after delay1 + 2850*delay_incr;
elsif nramp = '0' and StoredData = "101100100011" then SHout <= '1' after delay1 + 2851*delay_incr;
elsif nramp = '0' and StoredData = "101100100100" then SHout <= '1' after delay1 + 2852*delay_incr;
elsif nramp = '0' and StoredData = "101100100101" then SHout <= '1' after delay1 + 2853*delay_incr;
elsif nramp = '0' and StoredData = "101100100110" then SHout <= '1' after delay1 + 2854*delay_incr;
elsif nramp = '0' and StoredData = "101100100111" then SHout <= '1' after delay1 + 2855*delay_incr;
elsif nramp = '0' and StoredData = "101100101000" then SHout <= '1' after delay1 + 2856*delay_incr;
elsif nramp = '0' and StoredData = "101100101001" then SHout <= '1' after delay1 + 2857*delay_incr;
elsif nramp = '0' and StoredData = "101100101010" then SHout <= '1' after delay1 + 2858*delay_incr;
elsif nramp = '0' and StoredData = "101100101011" then SHout <= '1' after delay1 + 2859*delay_incr;
elsif nramp = '0' and StoredData = "101100101100" then SHout <= '1' after delay1 + 2860*delay_incr;
elsif nramp = '0' and StoredData = "101100101101" then SHout <= '1' after delay1 + 2861*delay_incr;
elsif nramp = '0' and StoredData = "101100101110" then SHout <= '1' after delay1 + 2862*delay_incr;
elsif nramp = '0' and StoredData = "101100101111" then SHout <= '1' after delay1 + 2863*delay_incr;
elsif nramp = '0' and StoredData = "101100110000" then SHout <= '1' after delay1 + 2864*delay_incr;
elsif nramp = '0' and StoredData = "101100110001" then SHout <= '1' after delay1 + 2865*delay_incr;
elsif nramp = '0' and StoredData = "101100110010" then SHout <= '1' after delay1 + 2866*delay_incr;
elsif nramp = '0' and StoredData = "101100110011" then SHout <= '1' after delay1 + 2867*delay_incr;
elsif nramp = '0' and StoredData = "101100110100" then SHout <= '1' after delay1 + 2868*delay_incr;
elsif nramp = '0' and StoredData = "101100110101" then SHout <= '1' after delay1 + 2869*delay_incr;
elsif nramp = '0' and StoredData = "101100110110" then SHout <= '1' after delay1 + 2870*delay_incr;
elsif nramp = '0' and StoredData = "101100110111" then SHout <= '1' after delay1 + 2871*delay_incr;
elsif nramp = '0' and StoredData = "101100111000" then SHout <= '1' after delay1 + 2872*delay_incr;
elsif nramp = '0' and StoredData = "101100111001" then SHout <= '1' after delay1 + 2873*delay_incr;
elsif nramp = '0' and StoredData = "101100111010" then SHout <= '1' after delay1 + 2874*delay_incr;
elsif nramp = '0' and StoredData = "101100111011" then SHout <= '1' after delay1 + 2875*delay_incr;
elsif nramp = '0' and StoredData = "101100111100" then SHout <= '1' after delay1 + 2876*delay_incr;
elsif nramp = '0' and StoredData = "101100111101" then SHout <= '1' after delay1 + 2877*delay_incr;
elsif nramp = '0' and StoredData = "101100111110" then SHout <= '1' after delay1 + 2878*delay_incr;
elsif nramp = '0' and StoredData = "101100111111" then SHout <= '1' after delay1 + 2879*delay_incr;
elsif nramp = '0' and StoredData = "101101000000" then SHout <= '1' after delay1 + 2880*delay_incr;
elsif nramp = '0' and StoredData = "101101000001" then SHout <= '1' after delay1 + 2881*delay_incr;
elsif nramp = '0' and StoredData = "101101000010" then SHout <= '1' after delay1 + 2882*delay_incr;
elsif nramp = '0' and StoredData = "101101000011" then SHout <= '1' after delay1 + 2883*delay_incr;
elsif nramp = '0' and StoredData = "101101000100" then SHout <= '1' after delay1 + 2884*delay_incr;
elsif nramp = '0' and StoredData = "101101000101" then SHout <= '1' after delay1 + 2885*delay_incr;
elsif nramp = '0' and StoredData = "101101000110" then SHout <= '1' after delay1 + 2886*delay_incr;
elsif nramp = '0' and StoredData = "101101000111" then SHout <= '1' after delay1 + 2887*delay_incr;
elsif nramp = '0' and StoredData = "101101001000" then SHout <= '1' after delay1 + 2888*delay_incr;
elsif nramp = '0' and StoredData = "101101001001" then SHout <= '1' after delay1 + 2889*delay_incr;
elsif nramp = '0' and StoredData = "101101001010" then SHout <= '1' after delay1 + 2890*delay_incr;
elsif nramp = '0' and StoredData = "101101001011" then SHout <= '1' after delay1 + 2891*delay_incr;
elsif nramp = '0' and StoredData = "101101001100" then SHout <= '1' after delay1 + 2892*delay_incr;
elsif nramp = '0' and StoredData = "101101001101" then SHout <= '1' after delay1 + 2893*delay_incr;
elsif nramp = '0' and StoredData = "101101001110" then SHout <= '1' after delay1 + 2894*delay_incr;
elsif nramp = '0' and StoredData = "101101001111" then SHout <= '1' after delay1 + 2895*delay_incr;
elsif nramp = '0' and StoredData = "101101010000" then SHout <= '1' after delay1 + 2896*delay_incr;
elsif nramp = '0' and StoredData = "101101010001" then SHout <= '1' after delay1 + 2897*delay_incr;
elsif nramp = '0' and StoredData = "101101010010" then SHout <= '1' after delay1 + 2898*delay_incr;
elsif nramp = '0' and StoredData = "101101010011" then SHout <= '1' after delay1 + 2899*delay_incr;
elsif nramp = '0' and StoredData = "101101010100" then SHout <= '1' after delay1 + 2900*delay_incr;
elsif nramp = '0' and StoredData = "101101010101" then SHout <= '1' after delay1 + 2901*delay_incr;
elsif nramp = '0' and StoredData = "101101010110" then SHout <= '1' after delay1 + 2902*delay_incr;
elsif nramp = '0' and StoredData = "101101010111" then SHout <= '1' after delay1 + 2903*delay_incr;
elsif nramp = '0' and StoredData = "101101011000" then SHout <= '1' after delay1 + 2904*delay_incr;
elsif nramp = '0' and StoredData = "101101011001" then SHout <= '1' after delay1 + 2905*delay_incr;
elsif nramp = '0' and StoredData = "101101011010" then SHout <= '1' after delay1 + 2906*delay_incr;
elsif nramp = '0' and StoredData = "101101011011" then SHout <= '1' after delay1 + 2907*delay_incr;
elsif nramp = '0' and StoredData = "101101011100" then SHout <= '1' after delay1 + 2908*delay_incr;
elsif nramp = '0' and StoredData = "101101011101" then SHout <= '1' after delay1 + 2909*delay_incr;
elsif nramp = '0' and StoredData = "101101011110" then SHout <= '1' after delay1 + 2910*delay_incr;
elsif nramp = '0' and StoredData = "101101011111" then SHout <= '1' after delay1 + 2911*delay_incr;
elsif nramp = '0' and StoredData = "101101100000" then SHout <= '1' after delay1 + 2912*delay_incr;
elsif nramp = '0' and StoredData = "101101100001" then SHout <= '1' after delay1 + 2913*delay_incr;
elsif nramp = '0' and StoredData = "101101100010" then SHout <= '1' after delay1 + 2914*delay_incr;
elsif nramp = '0' and StoredData = "101101100011" then SHout <= '1' after delay1 + 2915*delay_incr;
elsif nramp = '0' and StoredData = "101101100100" then SHout <= '1' after delay1 + 2916*delay_incr;
elsif nramp = '0' and StoredData = "101101100101" then SHout <= '1' after delay1 + 2917*delay_incr;
elsif nramp = '0' and StoredData = "101101100110" then SHout <= '1' after delay1 + 2918*delay_incr;
elsif nramp = '0' and StoredData = "101101100111" then SHout <= '1' after delay1 + 2919*delay_incr;
elsif nramp = '0' and StoredData = "101101101000" then SHout <= '1' after delay1 + 2920*delay_incr;
elsif nramp = '0' and StoredData = "101101101001" then SHout <= '1' after delay1 + 2921*delay_incr;
elsif nramp = '0' and StoredData = "101101101010" then SHout <= '1' after delay1 + 2922*delay_incr;
elsif nramp = '0' and StoredData = "101101101011" then SHout <= '1' after delay1 + 2923*delay_incr;
elsif nramp = '0' and StoredData = "101101101100" then SHout <= '1' after delay1 + 2924*delay_incr;
elsif nramp = '0' and StoredData = "101101101101" then SHout <= '1' after delay1 + 2925*delay_incr;
elsif nramp = '0' and StoredData = "101101101110" then SHout <= '1' after delay1 + 2926*delay_incr;
elsif nramp = '0' and StoredData = "101101101111" then SHout <= '1' after delay1 + 2927*delay_incr;
elsif nramp = '0' and StoredData = "101101110000" then SHout <= '1' after delay1 + 2928*delay_incr;
elsif nramp = '0' and StoredData = "101101110001" then SHout <= '1' after delay1 + 2929*delay_incr;
elsif nramp = '0' and StoredData = "101101110010" then SHout <= '1' after delay1 + 2930*delay_incr;
elsif nramp = '0' and StoredData = "101101110011" then SHout <= '1' after delay1 + 2931*delay_incr;
elsif nramp = '0' and StoredData = "101101110100" then SHout <= '1' after delay1 + 2932*delay_incr;
elsif nramp = '0' and StoredData = "101101110101" then SHout <= '1' after delay1 + 2933*delay_incr;
elsif nramp = '0' and StoredData = "101101110110" then SHout <= '1' after delay1 + 2934*delay_incr;
elsif nramp = '0' and StoredData = "101101110111" then SHout <= '1' after delay1 + 2935*delay_incr;
elsif nramp = '0' and StoredData = "101101111000" then SHout <= '1' after delay1 + 2936*delay_incr;
elsif nramp = '0' and StoredData = "101101111001" then SHout <= '1' after delay1 + 2937*delay_incr;
elsif nramp = '0' and StoredData = "101101111010" then SHout <= '1' after delay1 + 2938*delay_incr;
elsif nramp = '0' and StoredData = "101101111011" then SHout <= '1' after delay1 + 2939*delay_incr;
elsif nramp = '0' and StoredData = "101101111100" then SHout <= '1' after delay1 + 2940*delay_incr;
elsif nramp = '0' and StoredData = "101101111101" then SHout <= '1' after delay1 + 2941*delay_incr;
elsif nramp = '0' and StoredData = "101101111110" then SHout <= '1' after delay1 + 2942*delay_incr;
elsif nramp = '0' and StoredData = "101101111111" then SHout <= '1' after delay1 + 2943*delay_incr;
elsif nramp = '0' and StoredData = "101110000000" then SHout <= '1' after delay1 + 2944*delay_incr;
elsif nramp = '0' and StoredData = "101110000001" then SHout <= '1' after delay1 + 2945*delay_incr;
elsif nramp = '0' and StoredData = "101110000010" then SHout <= '1' after delay1 + 2946*delay_incr;
elsif nramp = '0' and StoredData = "101110000011" then SHout <= '1' after delay1 + 2947*delay_incr;
elsif nramp = '0' and StoredData = "101110000100" then SHout <= '1' after delay1 + 2948*delay_incr;
elsif nramp = '0' and StoredData = "101110000101" then SHout <= '1' after delay1 + 2949*delay_incr;
elsif nramp = '0' and StoredData = "101110000110" then SHout <= '1' after delay1 + 2950*delay_incr;
elsif nramp = '0' and StoredData = "101110000111" then SHout <= '1' after delay1 + 2951*delay_incr;
elsif nramp = '0' and StoredData = "101110001000" then SHout <= '1' after delay1 + 2952*delay_incr;
elsif nramp = '0' and StoredData = "101110001001" then SHout <= '1' after delay1 + 2953*delay_incr;
elsif nramp = '0' and StoredData = "101110001010" then SHout <= '1' after delay1 + 2954*delay_incr;
elsif nramp = '0' and StoredData = "101110001011" then SHout <= '1' after delay1 + 2955*delay_incr;
elsif nramp = '0' and StoredData = "101110001100" then SHout <= '1' after delay1 + 2956*delay_incr;
elsif nramp = '0' and StoredData = "101110001101" then SHout <= '1' after delay1 + 2957*delay_incr;
elsif nramp = '0' and StoredData = "101110001110" then SHout <= '1' after delay1 + 2958*delay_incr;
elsif nramp = '0' and StoredData = "101110001111" then SHout <= '1' after delay1 + 2959*delay_incr;
elsif nramp = '0' and StoredData = "101110010000" then SHout <= '1' after delay1 + 2960*delay_incr;
elsif nramp = '0' and StoredData = "101110010001" then SHout <= '1' after delay1 + 2961*delay_incr;
elsif nramp = '0' and StoredData = "101110010010" then SHout <= '1' after delay1 + 2962*delay_incr;
elsif nramp = '0' and StoredData = "101110010011" then SHout <= '1' after delay1 + 2963*delay_incr;
elsif nramp = '0' and StoredData = "101110010100" then SHout <= '1' after delay1 + 2964*delay_incr;
elsif nramp = '0' and StoredData = "101110010101" then SHout <= '1' after delay1 + 2965*delay_incr;
elsif nramp = '0' and StoredData = "101110010110" then SHout <= '1' after delay1 + 2966*delay_incr;
elsif nramp = '0' and StoredData = "101110010111" then SHout <= '1' after delay1 + 2967*delay_incr;
elsif nramp = '0' and StoredData = "101110011000" then SHout <= '1' after delay1 + 2968*delay_incr;
elsif nramp = '0' and StoredData = "101110011001" then SHout <= '1' after delay1 + 2969*delay_incr;
elsif nramp = '0' and StoredData = "101110011010" then SHout <= '1' after delay1 + 2970*delay_incr;
elsif nramp = '0' and StoredData = "101110011011" then SHout <= '1' after delay1 + 2971*delay_incr;
elsif nramp = '0' and StoredData = "101110011100" then SHout <= '1' after delay1 + 2972*delay_incr;
elsif nramp = '0' and StoredData = "101110011101" then SHout <= '1' after delay1 + 2973*delay_incr;
elsif nramp = '0' and StoredData = "101110011110" then SHout <= '1' after delay1 + 2974*delay_incr;
elsif nramp = '0' and StoredData = "101110011111" then SHout <= '1' after delay1 + 2975*delay_incr;
elsif nramp = '0' and StoredData = "101110100000" then SHout <= '1' after delay1 + 2976*delay_incr;
elsif nramp = '0' and StoredData = "101110100001" then SHout <= '1' after delay1 + 2977*delay_incr;
elsif nramp = '0' and StoredData = "101110100010" then SHout <= '1' after delay1 + 2978*delay_incr;
elsif nramp = '0' and StoredData = "101110100011" then SHout <= '1' after delay1 + 2979*delay_incr;
elsif nramp = '0' and StoredData = "101110100100" then SHout <= '1' after delay1 + 2980*delay_incr;
elsif nramp = '0' and StoredData = "101110100101" then SHout <= '1' after delay1 + 2981*delay_incr;
elsif nramp = '0' and StoredData = "101110100110" then SHout <= '1' after delay1 + 2982*delay_incr;
elsif nramp = '0' and StoredData = "101110100111" then SHout <= '1' after delay1 + 2983*delay_incr;
elsif nramp = '0' and StoredData = "101110101000" then SHout <= '1' after delay1 + 2984*delay_incr;
elsif nramp = '0' and StoredData = "101110101001" then SHout <= '1' after delay1 + 2985*delay_incr;
elsif nramp = '0' and StoredData = "101110101010" then SHout <= '1' after delay1 + 2986*delay_incr;
elsif nramp = '0' and StoredData = "101110101011" then SHout <= '1' after delay1 + 2987*delay_incr;
elsif nramp = '0' and StoredData = "101110101100" then SHout <= '1' after delay1 + 2988*delay_incr;
elsif nramp = '0' and StoredData = "101110101101" then SHout <= '1' after delay1 + 2989*delay_incr;
elsif nramp = '0' and StoredData = "101110101110" then SHout <= '1' after delay1 + 2990*delay_incr;
elsif nramp = '0' and StoredData = "101110101111" then SHout <= '1' after delay1 + 2991*delay_incr;
elsif nramp = '0' and StoredData = "101110110000" then SHout <= '1' after delay1 + 2992*delay_incr;
elsif nramp = '0' and StoredData = "101110110001" then SHout <= '1' after delay1 + 2993*delay_incr;
elsif nramp = '0' and StoredData = "101110110010" then SHout <= '1' after delay1 + 2994*delay_incr;
elsif nramp = '0' and StoredData = "101110110011" then SHout <= '1' after delay1 + 2995*delay_incr;
elsif nramp = '0' and StoredData = "101110110100" then SHout <= '1' after delay1 + 2996*delay_incr;
elsif nramp = '0' and StoredData = "101110110101" then SHout <= '1' after delay1 + 2997*delay_incr;
elsif nramp = '0' and StoredData = "101110110110" then SHout <= '1' after delay1 + 2998*delay_incr;
elsif nramp = '0' and StoredData = "101110110111" then SHout <= '1' after delay1 + 2999*delay_incr;
elsif nramp = '0' and StoredData = "101110111000" then SHout <= '1' after delay1 + 3000*delay_incr;
elsif nramp = '0' and StoredData = "101110111001" then SHout <= '1' after delay1 + 3001*delay_incr;
elsif nramp = '0' and StoredData = "101110111010" then SHout <= '1' after delay1 + 3002*delay_incr;
elsif nramp = '0' and StoredData = "101110111011" then SHout <= '1' after delay1 + 3003*delay_incr;
elsif nramp = '0' and StoredData = "101110111100" then SHout <= '1' after delay1 + 3004*delay_incr;
elsif nramp = '0' and StoredData = "101110111101" then SHout <= '1' after delay1 + 3005*delay_incr;
elsif nramp = '0' and StoredData = "101110111110" then SHout <= '1' after delay1 + 3006*delay_incr;
elsif nramp = '0' and StoredData = "101110111111" then SHout <= '1' after delay1 + 3007*delay_incr;
elsif nramp = '0' and StoredData = "101111000000" then SHout <= '1' after delay1 + 3008*delay_incr;
elsif nramp = '0' and StoredData = "101111000001" then SHout <= '1' after delay1 + 3009*delay_incr;
elsif nramp = '0' and StoredData = "101111000010" then SHout <= '1' after delay1 + 3010*delay_incr;
elsif nramp = '0' and StoredData = "101111000011" then SHout <= '1' after delay1 + 3011*delay_incr;
elsif nramp = '0' and StoredData = "101111000100" then SHout <= '1' after delay1 + 3012*delay_incr;
elsif nramp = '0' and StoredData = "101111000101" then SHout <= '1' after delay1 + 3013*delay_incr;
elsif nramp = '0' and StoredData = "101111000110" then SHout <= '1' after delay1 + 3014*delay_incr;
elsif nramp = '0' and StoredData = "101111000111" then SHout <= '1' after delay1 + 3015*delay_incr;
elsif nramp = '0' and StoredData = "101111001000" then SHout <= '1' after delay1 + 3016*delay_incr;
elsif nramp = '0' and StoredData = "101111001001" then SHout <= '1' after delay1 + 3017*delay_incr;
elsif nramp = '0' and StoredData = "101111001010" then SHout <= '1' after delay1 + 3018*delay_incr;
elsif nramp = '0' and StoredData = "101111001011" then SHout <= '1' after delay1 + 3019*delay_incr;
elsif nramp = '0' and StoredData = "101111001100" then SHout <= '1' after delay1 + 3020*delay_incr;
elsif nramp = '0' and StoredData = "101111001101" then SHout <= '1' after delay1 + 3021*delay_incr;
elsif nramp = '0' and StoredData = "101111001110" then SHout <= '1' after delay1 + 3022*delay_incr;
elsif nramp = '0' and StoredData = "101111001111" then SHout <= '1' after delay1 + 3023*delay_incr;
elsif nramp = '0' and StoredData = "101111010000" then SHout <= '1' after delay1 + 3024*delay_incr;
elsif nramp = '0' and StoredData = "101111010001" then SHout <= '1' after delay1 + 3025*delay_incr;
elsif nramp = '0' and StoredData = "101111010010" then SHout <= '1' after delay1 + 3026*delay_incr;
elsif nramp = '0' and StoredData = "101111010011" then SHout <= '1' after delay1 + 3027*delay_incr;
elsif nramp = '0' and StoredData = "101111010100" then SHout <= '1' after delay1 + 3028*delay_incr;
elsif nramp = '0' and StoredData = "101111010101" then SHout <= '1' after delay1 + 3029*delay_incr;
elsif nramp = '0' and StoredData = "101111010110" then SHout <= '1' after delay1 + 3030*delay_incr;
elsif nramp = '0' and StoredData = "101111010111" then SHout <= '1' after delay1 + 3031*delay_incr;
elsif nramp = '0' and StoredData = "101111011000" then SHout <= '1' after delay1 + 3032*delay_incr;
elsif nramp = '0' and StoredData = "101111011001" then SHout <= '1' after delay1 + 3033*delay_incr;
elsif nramp = '0' and StoredData = "101111011010" then SHout <= '1' after delay1 + 3034*delay_incr;
elsif nramp = '0' and StoredData = "101111011011" then SHout <= '1' after delay1 + 3035*delay_incr;
elsif nramp = '0' and StoredData = "101111011100" then SHout <= '1' after delay1 + 3036*delay_incr;
elsif nramp = '0' and StoredData = "101111011101" then SHout <= '1' after delay1 + 3037*delay_incr;
elsif nramp = '0' and StoredData = "101111011110" then SHout <= '1' after delay1 + 3038*delay_incr;
elsif nramp = '0' and StoredData = "101111011111" then SHout <= '1' after delay1 + 3039*delay_incr;
elsif nramp = '0' and StoredData = "101111100000" then SHout <= '1' after delay1 + 3040*delay_incr;
elsif nramp = '0' and StoredData = "101111100001" then SHout <= '1' after delay1 + 3041*delay_incr;
elsif nramp = '0' and StoredData = "101111100010" then SHout <= '1' after delay1 + 3042*delay_incr;
elsif nramp = '0' and StoredData = "101111100011" then SHout <= '1' after delay1 + 3043*delay_incr;
elsif nramp = '0' and StoredData = "101111100100" then SHout <= '1' after delay1 + 3044*delay_incr;
elsif nramp = '0' and StoredData = "101111100101" then SHout <= '1' after delay1 + 3045*delay_incr;
elsif nramp = '0' and StoredData = "101111100110" then SHout <= '1' after delay1 + 3046*delay_incr;
elsif nramp = '0' and StoredData = "101111100111" then SHout <= '1' after delay1 + 3047*delay_incr;
elsif nramp = '0' and StoredData = "101111101000" then SHout <= '1' after delay1 + 3048*delay_incr;
elsif nramp = '0' and StoredData = "101111101001" then SHout <= '1' after delay1 + 3049*delay_incr;
elsif nramp = '0' and StoredData = "101111101010" then SHout <= '1' after delay1 + 3050*delay_incr;
elsif nramp = '0' and StoredData = "101111101011" then SHout <= '1' after delay1 + 3051*delay_incr;
elsif nramp = '0' and StoredData = "101111101100" then SHout <= '1' after delay1 + 3052*delay_incr;
elsif nramp = '0' and StoredData = "101111101101" then SHout <= '1' after delay1 + 3053*delay_incr;
elsif nramp = '0' and StoredData = "101111101110" then SHout <= '1' after delay1 + 3054*delay_incr;
elsif nramp = '0' and StoredData = "101111101111" then SHout <= '1' after delay1 + 3055*delay_incr;
elsif nramp = '0' and StoredData = "101111110000" then SHout <= '1' after delay1 + 3056*delay_incr;
elsif nramp = '0' and StoredData = "101111110001" then SHout <= '1' after delay1 + 3057*delay_incr;
elsif nramp = '0' and StoredData = "101111110010" then SHout <= '1' after delay1 + 3058*delay_incr;
elsif nramp = '0' and StoredData = "101111110011" then SHout <= '1' after delay1 + 3059*delay_incr;
elsif nramp = '0' and StoredData = "101111110100" then SHout <= '1' after delay1 + 3060*delay_incr;
elsif nramp = '0' and StoredData = "101111110101" then SHout <= '1' after delay1 + 3061*delay_incr;
elsif nramp = '0' and StoredData = "101111110110" then SHout <= '1' after delay1 + 3062*delay_incr;
elsif nramp = '0' and StoredData = "101111110111" then SHout <= '1' after delay1 + 3063*delay_incr;
elsif nramp = '0' and StoredData = "101111111000" then SHout <= '1' after delay1 + 3064*delay_incr;
elsif nramp = '0' and StoredData = "101111111001" then SHout <= '1' after delay1 + 3065*delay_incr;
elsif nramp = '0' and StoredData = "101111111010" then SHout <= '1' after delay1 + 3066*delay_incr;
elsif nramp = '0' and StoredData = "101111111011" then SHout <= '1' after delay1 + 3067*delay_incr;
elsif nramp = '0' and StoredData = "101111111100" then SHout <= '1' after delay1 + 3068*delay_incr;
elsif nramp = '0' and StoredData = "101111111101" then SHout <= '1' after delay1 + 3069*delay_incr;
elsif nramp = '0' and StoredData = "101111111110" then SHout <= '1' after delay1 + 3070*delay_incr;
elsif nramp = '0' and StoredData = "101111111111" then SHout <= '1' after delay1 + 3071*delay_incr;
elsif nramp = '0' and StoredData = "110000000000" then SHout <= '1' after delay1 + 3072*delay_incr;
elsif nramp = '0' and StoredData = "110000000001" then SHout <= '1' after delay1 + 3073*delay_incr;
elsif nramp = '0' and StoredData = "110000000010" then SHout <= '1' after delay1 + 3074*delay_incr;
elsif nramp = '0' and StoredData = "110000000011" then SHout <= '1' after delay1 + 3075*delay_incr;
elsif nramp = '0' and StoredData = "110000000100" then SHout <= '1' after delay1 + 3076*delay_incr;
elsif nramp = '0' and StoredData = "110000000101" then SHout <= '1' after delay1 + 3077*delay_incr;
elsif nramp = '0' and StoredData = "110000000110" then SHout <= '1' after delay1 + 3078*delay_incr;
elsif nramp = '0' and StoredData = "110000000111" then SHout <= '1' after delay1 + 3079*delay_incr;
elsif nramp = '0' and StoredData = "110000001000" then SHout <= '1' after delay1 + 3080*delay_incr;
elsif nramp = '0' and StoredData = "110000001001" then SHout <= '1' after delay1 + 3081*delay_incr;
elsif nramp = '0' and StoredData = "110000001010" then SHout <= '1' after delay1 + 3082*delay_incr;
elsif nramp = '0' and StoredData = "110000001011" then SHout <= '1' after delay1 + 3083*delay_incr;
elsif nramp = '0' and StoredData = "110000001100" then SHout <= '1' after delay1 + 3084*delay_incr;
elsif nramp = '0' and StoredData = "110000001101" then SHout <= '1' after delay1 + 3085*delay_incr;
elsif nramp = '0' and StoredData = "110000001110" then SHout <= '1' after delay1 + 3086*delay_incr;
elsif nramp = '0' and StoredData = "110000001111" then SHout <= '1' after delay1 + 3087*delay_incr;
elsif nramp = '0' and StoredData = "110000010000" then SHout <= '1' after delay1 + 3088*delay_incr;
elsif nramp = '0' and StoredData = "110000010001" then SHout <= '1' after delay1 + 3089*delay_incr;
elsif nramp = '0' and StoredData = "110000010010" then SHout <= '1' after delay1 + 3090*delay_incr;
elsif nramp = '0' and StoredData = "110000010011" then SHout <= '1' after delay1 + 3091*delay_incr;
elsif nramp = '0' and StoredData = "110000010100" then SHout <= '1' after delay1 + 3092*delay_incr;
elsif nramp = '0' and StoredData = "110000010101" then SHout <= '1' after delay1 + 3093*delay_incr;
elsif nramp = '0' and StoredData = "110000010110" then SHout <= '1' after delay1 + 3094*delay_incr;
elsif nramp = '0' and StoredData = "110000010111" then SHout <= '1' after delay1 + 3095*delay_incr;
elsif nramp = '0' and StoredData = "110000011000" then SHout <= '1' after delay1 + 3096*delay_incr;
elsif nramp = '0' and StoredData = "110000011001" then SHout <= '1' after delay1 + 3097*delay_incr;
elsif nramp = '0' and StoredData = "110000011010" then SHout <= '1' after delay1 + 3098*delay_incr;
elsif nramp = '0' and StoredData = "110000011011" then SHout <= '1' after delay1 + 3099*delay_incr;
elsif nramp = '0' and StoredData = "110000011100" then SHout <= '1' after delay1 + 3100*delay_incr;
elsif nramp = '0' and StoredData = "110000011101" then SHout <= '1' after delay1 + 3101*delay_incr;
elsif nramp = '0' and StoredData = "110000011110" then SHout <= '1' after delay1 + 3102*delay_incr;
elsif nramp = '0' and StoredData = "110000011111" then SHout <= '1' after delay1 + 3103*delay_incr;
elsif nramp = '0' and StoredData = "110000100000" then SHout <= '1' after delay1 + 3104*delay_incr;
elsif nramp = '0' and StoredData = "110000100001" then SHout <= '1' after delay1 + 3105*delay_incr;
elsif nramp = '0' and StoredData = "110000100010" then SHout <= '1' after delay1 + 3106*delay_incr;
elsif nramp = '0' and StoredData = "110000100011" then SHout <= '1' after delay1 + 3107*delay_incr;
elsif nramp = '0' and StoredData = "110000100100" then SHout <= '1' after delay1 + 3108*delay_incr;
elsif nramp = '0' and StoredData = "110000100101" then SHout <= '1' after delay1 + 3109*delay_incr;
elsif nramp = '0' and StoredData = "110000100110" then SHout <= '1' after delay1 + 3110*delay_incr;
elsif nramp = '0' and StoredData = "110000100111" then SHout <= '1' after delay1 + 3111*delay_incr;
elsif nramp = '0' and StoredData = "110000101000" then SHout <= '1' after delay1 + 3112*delay_incr;
elsif nramp = '0' and StoredData = "110000101001" then SHout <= '1' after delay1 + 3113*delay_incr;
elsif nramp = '0' and StoredData = "110000101010" then SHout <= '1' after delay1 + 3114*delay_incr;
elsif nramp = '0' and StoredData = "110000101011" then SHout <= '1' after delay1 + 3115*delay_incr;
elsif nramp = '0' and StoredData = "110000101100" then SHout <= '1' after delay1 + 3116*delay_incr;
elsif nramp = '0' and StoredData = "110000101101" then SHout <= '1' after delay1 + 3117*delay_incr;
elsif nramp = '0' and StoredData = "110000101110" then SHout <= '1' after delay1 + 3118*delay_incr;
elsif nramp = '0' and StoredData = "110000101111" then SHout <= '1' after delay1 + 3119*delay_incr;
elsif nramp = '0' and StoredData = "110000110000" then SHout <= '1' after delay1 + 3120*delay_incr;
elsif nramp = '0' and StoredData = "110000110001" then SHout <= '1' after delay1 + 3121*delay_incr;
elsif nramp = '0' and StoredData = "110000110010" then SHout <= '1' after delay1 + 3122*delay_incr;
elsif nramp = '0' and StoredData = "110000110011" then SHout <= '1' after delay1 + 3123*delay_incr;
elsif nramp = '0' and StoredData = "110000110100" then SHout <= '1' after delay1 + 3124*delay_incr;
elsif nramp = '0' and StoredData = "110000110101" then SHout <= '1' after delay1 + 3125*delay_incr;
elsif nramp = '0' and StoredData = "110000110110" then SHout <= '1' after delay1 + 3126*delay_incr;
elsif nramp = '0' and StoredData = "110000110111" then SHout <= '1' after delay1 + 3127*delay_incr;
elsif nramp = '0' and StoredData = "110000111000" then SHout <= '1' after delay1 + 3128*delay_incr;
elsif nramp = '0' and StoredData = "110000111001" then SHout <= '1' after delay1 + 3129*delay_incr;
elsif nramp = '0' and StoredData = "110000111010" then SHout <= '1' after delay1 + 3130*delay_incr;
elsif nramp = '0' and StoredData = "110000111011" then SHout <= '1' after delay1 + 3131*delay_incr;
elsif nramp = '0' and StoredData = "110000111100" then SHout <= '1' after delay1 + 3132*delay_incr;
elsif nramp = '0' and StoredData = "110000111101" then SHout <= '1' after delay1 + 3133*delay_incr;
elsif nramp = '0' and StoredData = "110000111110" then SHout <= '1' after delay1 + 3134*delay_incr;
elsif nramp = '0' and StoredData = "110000111111" then SHout <= '1' after delay1 + 3135*delay_incr;
elsif nramp = '0' and StoredData = "110001000000" then SHout <= '1' after delay1 + 3136*delay_incr;
elsif nramp = '0' and StoredData = "110001000001" then SHout <= '1' after delay1 + 3137*delay_incr;
elsif nramp = '0' and StoredData = "110001000010" then SHout <= '1' after delay1 + 3138*delay_incr;
elsif nramp = '0' and StoredData = "110001000011" then SHout <= '1' after delay1 + 3139*delay_incr;
elsif nramp = '0' and StoredData = "110001000100" then SHout <= '1' after delay1 + 3140*delay_incr;
elsif nramp = '0' and StoredData = "110001000101" then SHout <= '1' after delay1 + 3141*delay_incr;
elsif nramp = '0' and StoredData = "110001000110" then SHout <= '1' after delay1 + 3142*delay_incr;
elsif nramp = '0' and StoredData = "110001000111" then SHout <= '1' after delay1 + 3143*delay_incr;
elsif nramp = '0' and StoredData = "110001001000" then SHout <= '1' after delay1 + 3144*delay_incr;
elsif nramp = '0' and StoredData = "110001001001" then SHout <= '1' after delay1 + 3145*delay_incr;
elsif nramp = '0' and StoredData = "110001001010" then SHout <= '1' after delay1 + 3146*delay_incr;
elsif nramp = '0' and StoredData = "110001001011" then SHout <= '1' after delay1 + 3147*delay_incr;
elsif nramp = '0' and StoredData = "110001001100" then SHout <= '1' after delay1 + 3148*delay_incr;
elsif nramp = '0' and StoredData = "110001001101" then SHout <= '1' after delay1 + 3149*delay_incr;
elsif nramp = '0' and StoredData = "110001001110" then SHout <= '1' after delay1 + 3150*delay_incr;
elsif nramp = '0' and StoredData = "110001001111" then SHout <= '1' after delay1 + 3151*delay_incr;
elsif nramp = '0' and StoredData = "110001010000" then SHout <= '1' after delay1 + 3152*delay_incr;
elsif nramp = '0' and StoredData = "110001010001" then SHout <= '1' after delay1 + 3153*delay_incr;
elsif nramp = '0' and StoredData = "110001010010" then SHout <= '1' after delay1 + 3154*delay_incr;
elsif nramp = '0' and StoredData = "110001010011" then SHout <= '1' after delay1 + 3155*delay_incr;
elsif nramp = '0' and StoredData = "110001010100" then SHout <= '1' after delay1 + 3156*delay_incr;
elsif nramp = '0' and StoredData = "110001010101" then SHout <= '1' after delay1 + 3157*delay_incr;
elsif nramp = '0' and StoredData = "110001010110" then SHout <= '1' after delay1 + 3158*delay_incr;
elsif nramp = '0' and StoredData = "110001010111" then SHout <= '1' after delay1 + 3159*delay_incr;
elsif nramp = '0' and StoredData = "110001011000" then SHout <= '1' after delay1 + 3160*delay_incr;
elsif nramp = '0' and StoredData = "110001011001" then SHout <= '1' after delay1 + 3161*delay_incr;
elsif nramp = '0' and StoredData = "110001011010" then SHout <= '1' after delay1 + 3162*delay_incr;
elsif nramp = '0' and StoredData = "110001011011" then SHout <= '1' after delay1 + 3163*delay_incr;
elsif nramp = '0' and StoredData = "110001011100" then SHout <= '1' after delay1 + 3164*delay_incr;
elsif nramp = '0' and StoredData = "110001011101" then SHout <= '1' after delay1 + 3165*delay_incr;
elsif nramp = '0' and StoredData = "110001011110" then SHout <= '1' after delay1 + 3166*delay_incr;
elsif nramp = '0' and StoredData = "110001011111" then SHout <= '1' after delay1 + 3167*delay_incr;
elsif nramp = '0' and StoredData = "110001100000" then SHout <= '1' after delay1 + 3168*delay_incr;
elsif nramp = '0' and StoredData = "110001100001" then SHout <= '1' after delay1 + 3169*delay_incr;
elsif nramp = '0' and StoredData = "110001100010" then SHout <= '1' after delay1 + 3170*delay_incr;
elsif nramp = '0' and StoredData = "110001100011" then SHout <= '1' after delay1 + 3171*delay_incr;
elsif nramp = '0' and StoredData = "110001100100" then SHout <= '1' after delay1 + 3172*delay_incr;
elsif nramp = '0' and StoredData = "110001100101" then SHout <= '1' after delay1 + 3173*delay_incr;
elsif nramp = '0' and StoredData = "110001100110" then SHout <= '1' after delay1 + 3174*delay_incr;
elsif nramp = '0' and StoredData = "110001100111" then SHout <= '1' after delay1 + 3175*delay_incr;
elsif nramp = '0' and StoredData = "110001101000" then SHout <= '1' after delay1 + 3176*delay_incr;
elsif nramp = '0' and StoredData = "110001101001" then SHout <= '1' after delay1 + 3177*delay_incr;
elsif nramp = '0' and StoredData = "110001101010" then SHout <= '1' after delay1 + 3178*delay_incr;
elsif nramp = '0' and StoredData = "110001101011" then SHout <= '1' after delay1 + 3179*delay_incr;
elsif nramp = '0' and StoredData = "110001101100" then SHout <= '1' after delay1 + 3180*delay_incr;
elsif nramp = '0' and StoredData = "110001101101" then SHout <= '1' after delay1 + 3181*delay_incr;
elsif nramp = '0' and StoredData = "110001101110" then SHout <= '1' after delay1 + 3182*delay_incr;
elsif nramp = '0' and StoredData = "110001101111" then SHout <= '1' after delay1 + 3183*delay_incr;
elsif nramp = '0' and StoredData = "110001110000" then SHout <= '1' after delay1 + 3184*delay_incr;
elsif nramp = '0' and StoredData = "110001110001" then SHout <= '1' after delay1 + 3185*delay_incr;
elsif nramp = '0' and StoredData = "110001110010" then SHout <= '1' after delay1 + 3186*delay_incr;
elsif nramp = '0' and StoredData = "110001110011" then SHout <= '1' after delay1 + 3187*delay_incr;
elsif nramp = '0' and StoredData = "110001110100" then SHout <= '1' after delay1 + 3188*delay_incr;
elsif nramp = '0' and StoredData = "110001110101" then SHout <= '1' after delay1 + 3189*delay_incr;
elsif nramp = '0' and StoredData = "110001110110" then SHout <= '1' after delay1 + 3190*delay_incr;
elsif nramp = '0' and StoredData = "110001110111" then SHout <= '1' after delay1 + 3191*delay_incr;
elsif nramp = '0' and StoredData = "110001111000" then SHout <= '1' after delay1 + 3192*delay_incr;
elsif nramp = '0' and StoredData = "110001111001" then SHout <= '1' after delay1 + 3193*delay_incr;
elsif nramp = '0' and StoredData = "110001111010" then SHout <= '1' after delay1 + 3194*delay_incr;
elsif nramp = '0' and StoredData = "110001111011" then SHout <= '1' after delay1 + 3195*delay_incr;
elsif nramp = '0' and StoredData = "110001111100" then SHout <= '1' after delay1 + 3196*delay_incr;
elsif nramp = '0' and StoredData = "110001111101" then SHout <= '1' after delay1 + 3197*delay_incr;
elsif nramp = '0' and StoredData = "110001111110" then SHout <= '1' after delay1 + 3198*delay_incr;
elsif nramp = '0' and StoredData = "110001111111" then SHout <= '1' after delay1 + 3199*delay_incr;
elsif nramp = '0' and StoredData = "110010000000" then SHout <= '1' after delay1 + 3200*delay_incr;
elsif nramp = '0' and StoredData = "110010000001" then SHout <= '1' after delay1 + 3201*delay_incr;
elsif nramp = '0' and StoredData = "110010000010" then SHout <= '1' after delay1 + 3202*delay_incr;
elsif nramp = '0' and StoredData = "110010000011" then SHout <= '1' after delay1 + 3203*delay_incr;
elsif nramp = '0' and StoredData = "110010000100" then SHout <= '1' after delay1 + 3204*delay_incr;
elsif nramp = '0' and StoredData = "110010000101" then SHout <= '1' after delay1 + 3205*delay_incr;
elsif nramp = '0' and StoredData = "110010000110" then SHout <= '1' after delay1 + 3206*delay_incr;
elsif nramp = '0' and StoredData = "110010000111" then SHout <= '1' after delay1 + 3207*delay_incr;
elsif nramp = '0' and StoredData = "110010001000" then SHout <= '1' after delay1 + 3208*delay_incr;
elsif nramp = '0' and StoredData = "110010001001" then SHout <= '1' after delay1 + 3209*delay_incr;
elsif nramp = '0' and StoredData = "110010001010" then SHout <= '1' after delay1 + 3210*delay_incr;
elsif nramp = '0' and StoredData = "110010001011" then SHout <= '1' after delay1 + 3211*delay_incr;
elsif nramp = '0' and StoredData = "110010001100" then SHout <= '1' after delay1 + 3212*delay_incr;
elsif nramp = '0' and StoredData = "110010001101" then SHout <= '1' after delay1 + 3213*delay_incr;
elsif nramp = '0' and StoredData = "110010001110" then SHout <= '1' after delay1 + 3214*delay_incr;
elsif nramp = '0' and StoredData = "110010001111" then SHout <= '1' after delay1 + 3215*delay_incr;
elsif nramp = '0' and StoredData = "110010010000" then SHout <= '1' after delay1 + 3216*delay_incr;
elsif nramp = '0' and StoredData = "110010010001" then SHout <= '1' after delay1 + 3217*delay_incr;
elsif nramp = '0' and StoredData = "110010010010" then SHout <= '1' after delay1 + 3218*delay_incr;
elsif nramp = '0' and StoredData = "110010010011" then SHout <= '1' after delay1 + 3219*delay_incr;
elsif nramp = '0' and StoredData = "110010010100" then SHout <= '1' after delay1 + 3220*delay_incr;
elsif nramp = '0' and StoredData = "110010010101" then SHout <= '1' after delay1 + 3221*delay_incr;
elsif nramp = '0' and StoredData = "110010010110" then SHout <= '1' after delay1 + 3222*delay_incr;
elsif nramp = '0' and StoredData = "110010010111" then SHout <= '1' after delay1 + 3223*delay_incr;
elsif nramp = '0' and StoredData = "110010011000" then SHout <= '1' after delay1 + 3224*delay_incr;
elsif nramp = '0' and StoredData = "110010011001" then SHout <= '1' after delay1 + 3225*delay_incr;
elsif nramp = '0' and StoredData = "110010011010" then SHout <= '1' after delay1 + 3226*delay_incr;
elsif nramp = '0' and StoredData = "110010011011" then SHout <= '1' after delay1 + 3227*delay_incr;
elsif nramp = '0' and StoredData = "110010011100" then SHout <= '1' after delay1 + 3228*delay_incr;
elsif nramp = '0' and StoredData = "110010011101" then SHout <= '1' after delay1 + 3229*delay_incr;
elsif nramp = '0' and StoredData = "110010011110" then SHout <= '1' after delay1 + 3230*delay_incr;
elsif nramp = '0' and StoredData = "110010011111" then SHout <= '1' after delay1 + 3231*delay_incr;
elsif nramp = '0' and StoredData = "110010100000" then SHout <= '1' after delay1 + 3232*delay_incr;
elsif nramp = '0' and StoredData = "110010100001" then SHout <= '1' after delay1 + 3233*delay_incr;
elsif nramp = '0' and StoredData = "110010100010" then SHout <= '1' after delay1 + 3234*delay_incr;
elsif nramp = '0' and StoredData = "110010100011" then SHout <= '1' after delay1 + 3235*delay_incr;
elsif nramp = '0' and StoredData = "110010100100" then SHout <= '1' after delay1 + 3236*delay_incr;
elsif nramp = '0' and StoredData = "110010100101" then SHout <= '1' after delay1 + 3237*delay_incr;
elsif nramp = '0' and StoredData = "110010100110" then SHout <= '1' after delay1 + 3238*delay_incr;
elsif nramp = '0' and StoredData = "110010100111" then SHout <= '1' after delay1 + 3239*delay_incr;
elsif nramp = '0' and StoredData = "110010101000" then SHout <= '1' after delay1 + 3240*delay_incr;
elsif nramp = '0' and StoredData = "110010101001" then SHout <= '1' after delay1 + 3241*delay_incr;
elsif nramp = '0' and StoredData = "110010101010" then SHout <= '1' after delay1 + 3242*delay_incr;
elsif nramp = '0' and StoredData = "110010101011" then SHout <= '1' after delay1 + 3243*delay_incr;
elsif nramp = '0' and StoredData = "110010101100" then SHout <= '1' after delay1 + 3244*delay_incr;
elsif nramp = '0' and StoredData = "110010101101" then SHout <= '1' after delay1 + 3245*delay_incr;
elsif nramp = '0' and StoredData = "110010101110" then SHout <= '1' after delay1 + 3246*delay_incr;
elsif nramp = '0' and StoredData = "110010101111" then SHout <= '1' after delay1 + 3247*delay_incr;
elsif nramp = '0' and StoredData = "110010110000" then SHout <= '1' after delay1 + 3248*delay_incr;
elsif nramp = '0' and StoredData = "110010110001" then SHout <= '1' after delay1 + 3249*delay_incr;
elsif nramp = '0' and StoredData = "110010110010" then SHout <= '1' after delay1 + 3250*delay_incr;
elsif nramp = '0' and StoredData = "110010110011" then SHout <= '1' after delay1 + 3251*delay_incr;
elsif nramp = '0' and StoredData = "110010110100" then SHout <= '1' after delay1 + 3252*delay_incr;
elsif nramp = '0' and StoredData = "110010110101" then SHout <= '1' after delay1 + 3253*delay_incr;
elsif nramp = '0' and StoredData = "110010110110" then SHout <= '1' after delay1 + 3254*delay_incr;
elsif nramp = '0' and StoredData = "110010110111" then SHout <= '1' after delay1 + 3255*delay_incr;
elsif nramp = '0' and StoredData = "110010111000" then SHout <= '1' after delay1 + 3256*delay_incr;
elsif nramp = '0' and StoredData = "110010111001" then SHout <= '1' after delay1 + 3257*delay_incr;
elsif nramp = '0' and StoredData = "110010111010" then SHout <= '1' after delay1 + 3258*delay_incr;
elsif nramp = '0' and StoredData = "110010111011" then SHout <= '1' after delay1 + 3259*delay_incr;
elsif nramp = '0' and StoredData = "110010111100" then SHout <= '1' after delay1 + 3260*delay_incr;
elsif nramp = '0' and StoredData = "110010111101" then SHout <= '1' after delay1 + 3261*delay_incr;
elsif nramp = '0' and StoredData = "110010111110" then SHout <= '1' after delay1 + 3262*delay_incr;
elsif nramp = '0' and StoredData = "110010111111" then SHout <= '1' after delay1 + 3263*delay_incr;
elsif nramp = '0' and StoredData = "110011000000" then SHout <= '1' after delay1 + 3264*delay_incr;
elsif nramp = '0' and StoredData = "110011000001" then SHout <= '1' after delay1 + 3265*delay_incr;
elsif nramp = '0' and StoredData = "110011000010" then SHout <= '1' after delay1 + 3266*delay_incr;
elsif nramp = '0' and StoredData = "110011000011" then SHout <= '1' after delay1 + 3267*delay_incr;
elsif nramp = '0' and StoredData = "110011000100" then SHout <= '1' after delay1 + 3268*delay_incr;
elsif nramp = '0' and StoredData = "110011000101" then SHout <= '1' after delay1 + 3269*delay_incr;
elsif nramp = '0' and StoredData = "110011000110" then SHout <= '1' after delay1 + 3270*delay_incr;
elsif nramp = '0' and StoredData = "110011000111" then SHout <= '1' after delay1 + 3271*delay_incr;
elsif nramp = '0' and StoredData = "110011001000" then SHout <= '1' after delay1 + 3272*delay_incr;
elsif nramp = '0' and StoredData = "110011001001" then SHout <= '1' after delay1 + 3273*delay_incr;
elsif nramp = '0' and StoredData = "110011001010" then SHout <= '1' after delay1 + 3274*delay_incr;
elsif nramp = '0' and StoredData = "110011001011" then SHout <= '1' after delay1 + 3275*delay_incr;
elsif nramp = '0' and StoredData = "110011001100" then SHout <= '1' after delay1 + 3276*delay_incr;
elsif nramp = '0' and StoredData = "110011001101" then SHout <= '1' after delay1 + 3277*delay_incr;
elsif nramp = '0' and StoredData = "110011001110" then SHout <= '1' after delay1 + 3278*delay_incr;
elsif nramp = '0' and StoredData = "110011001111" then SHout <= '1' after delay1 + 3279*delay_incr;
elsif nramp = '0' and StoredData = "110011010000" then SHout <= '1' after delay1 + 3280*delay_incr;
elsif nramp = '0' and StoredData = "110011010001" then SHout <= '1' after delay1 + 3281*delay_incr;
elsif nramp = '0' and StoredData = "110011010010" then SHout <= '1' after delay1 + 3282*delay_incr;
elsif nramp = '0' and StoredData = "110011010011" then SHout <= '1' after delay1 + 3283*delay_incr;
elsif nramp = '0' and StoredData = "110011010100" then SHout <= '1' after delay1 + 3284*delay_incr;
elsif nramp = '0' and StoredData = "110011010101" then SHout <= '1' after delay1 + 3285*delay_incr;
elsif nramp = '0' and StoredData = "110011010110" then SHout <= '1' after delay1 + 3286*delay_incr;
elsif nramp = '0' and StoredData = "110011010111" then SHout <= '1' after delay1 + 3287*delay_incr;
elsif nramp = '0' and StoredData = "110011011000" then SHout <= '1' after delay1 + 3288*delay_incr;
elsif nramp = '0' and StoredData = "110011011001" then SHout <= '1' after delay1 + 3289*delay_incr;
elsif nramp = '0' and StoredData = "110011011010" then SHout <= '1' after delay1 + 3290*delay_incr;
elsif nramp = '0' and StoredData = "110011011011" then SHout <= '1' after delay1 + 3291*delay_incr;
elsif nramp = '0' and StoredData = "110011011100" then SHout <= '1' after delay1 + 3292*delay_incr;
elsif nramp = '0' and StoredData = "110011011101" then SHout <= '1' after delay1 + 3293*delay_incr;
elsif nramp = '0' and StoredData = "110011011110" then SHout <= '1' after delay1 + 3294*delay_incr;
elsif nramp = '0' and StoredData = "110011011111" then SHout <= '1' after delay1 + 3295*delay_incr;
elsif nramp = '0' and StoredData = "110011100000" then SHout <= '1' after delay1 + 3296*delay_incr;
elsif nramp = '0' and StoredData = "110011100001" then SHout <= '1' after delay1 + 3297*delay_incr;
elsif nramp = '0' and StoredData = "110011100010" then SHout <= '1' after delay1 + 3298*delay_incr;
elsif nramp = '0' and StoredData = "110011100011" then SHout <= '1' after delay1 + 3299*delay_incr;
elsif nramp = '0' and StoredData = "110011100100" then SHout <= '1' after delay1 + 3300*delay_incr;
elsif nramp = '0' and StoredData = "110011100101" then SHout <= '1' after delay1 + 3301*delay_incr;
elsif nramp = '0' and StoredData = "110011100110" then SHout <= '1' after delay1 + 3302*delay_incr;
elsif nramp = '0' and StoredData = "110011100111" then SHout <= '1' after delay1 + 3303*delay_incr;
elsif nramp = '0' and StoredData = "110011101000" then SHout <= '1' after delay1 + 3304*delay_incr;
elsif nramp = '0' and StoredData = "110011101001" then SHout <= '1' after delay1 + 3305*delay_incr;
elsif nramp = '0' and StoredData = "110011101010" then SHout <= '1' after delay1 + 3306*delay_incr;
elsif nramp = '0' and StoredData = "110011101011" then SHout <= '1' after delay1 + 3307*delay_incr;
elsif nramp = '0' and StoredData = "110011101100" then SHout <= '1' after delay1 + 3308*delay_incr;
elsif nramp = '0' and StoredData = "110011101101" then SHout <= '1' after delay1 + 3309*delay_incr;
elsif nramp = '0' and StoredData = "110011101110" then SHout <= '1' after delay1 + 3310*delay_incr;
elsif nramp = '0' and StoredData = "110011101111" then SHout <= '1' after delay1 + 3311*delay_incr;
elsif nramp = '0' and StoredData = "110011110000" then SHout <= '1' after delay1 + 3312*delay_incr;
elsif nramp = '0' and StoredData = "110011110001" then SHout <= '1' after delay1 + 3313*delay_incr;
elsif nramp = '0' and StoredData = "110011110010" then SHout <= '1' after delay1 + 3314*delay_incr;
elsif nramp = '0' and StoredData = "110011110011" then SHout <= '1' after delay1 + 3315*delay_incr;
elsif nramp = '0' and StoredData = "110011110100" then SHout <= '1' after delay1 + 3316*delay_incr;
elsif nramp = '0' and StoredData = "110011110101" then SHout <= '1' after delay1 + 3317*delay_incr;
elsif nramp = '0' and StoredData = "110011110110" then SHout <= '1' after delay1 + 3318*delay_incr;
elsif nramp = '0' and StoredData = "110011110111" then SHout <= '1' after delay1 + 3319*delay_incr;
elsif nramp = '0' and StoredData = "110011111000" then SHout <= '1' after delay1 + 3320*delay_incr;
elsif nramp = '0' and StoredData = "110011111001" then SHout <= '1' after delay1 + 3321*delay_incr;
elsif nramp = '0' and StoredData = "110011111010" then SHout <= '1' after delay1 + 3322*delay_incr;
elsif nramp = '0' and StoredData = "110011111011" then SHout <= '1' after delay1 + 3323*delay_incr;
elsif nramp = '0' and StoredData = "110011111100" then SHout <= '1' after delay1 + 3324*delay_incr;
elsif nramp = '0' and StoredData = "110011111101" then SHout <= '1' after delay1 + 3325*delay_incr;
elsif nramp = '0' and StoredData = "110011111110" then SHout <= '1' after delay1 + 3326*delay_incr;
elsif nramp = '0' and StoredData = "110011111111" then SHout <= '1' after delay1 + 3327*delay_incr;
elsif nramp = '0' and StoredData = "110100000000" then SHout <= '1' after delay1 + 3328*delay_incr;
elsif nramp = '0' and StoredData = "110100000001" then SHout <= '1' after delay1 + 3329*delay_incr;
elsif nramp = '0' and StoredData = "110100000010" then SHout <= '1' after delay1 + 3330*delay_incr;
elsif nramp = '0' and StoredData = "110100000011" then SHout <= '1' after delay1 + 3331*delay_incr;
elsif nramp = '0' and StoredData = "110100000100" then SHout <= '1' after delay1 + 3332*delay_incr;
elsif nramp = '0' and StoredData = "110100000101" then SHout <= '1' after delay1 + 3333*delay_incr;
elsif nramp = '0' and StoredData = "110100000110" then SHout <= '1' after delay1 + 3334*delay_incr;
elsif nramp = '0' and StoredData = "110100000111" then SHout <= '1' after delay1 + 3335*delay_incr;
elsif nramp = '0' and StoredData = "110100001000" then SHout <= '1' after delay1 + 3336*delay_incr;
elsif nramp = '0' and StoredData = "110100001001" then SHout <= '1' after delay1 + 3337*delay_incr;
elsif nramp = '0' and StoredData = "110100001010" then SHout <= '1' after delay1 + 3338*delay_incr;
elsif nramp = '0' and StoredData = "110100001011" then SHout <= '1' after delay1 + 3339*delay_incr;
elsif nramp = '0' and StoredData = "110100001100" then SHout <= '1' after delay1 + 3340*delay_incr;
elsif nramp = '0' and StoredData = "110100001101" then SHout <= '1' after delay1 + 3341*delay_incr;
elsif nramp = '0' and StoredData = "110100001110" then SHout <= '1' after delay1 + 3342*delay_incr;
elsif nramp = '0' and StoredData = "110100001111" then SHout <= '1' after delay1 + 3343*delay_incr;
elsif nramp = '0' and StoredData = "110100010000" then SHout <= '1' after delay1 + 3344*delay_incr;
elsif nramp = '0' and StoredData = "110100010001" then SHout <= '1' after delay1 + 3345*delay_incr;
elsif nramp = '0' and StoredData = "110100010010" then SHout <= '1' after delay1 + 3346*delay_incr;
elsif nramp = '0' and StoredData = "110100010011" then SHout <= '1' after delay1 + 3347*delay_incr;
elsif nramp = '0' and StoredData = "110100010100" then SHout <= '1' after delay1 + 3348*delay_incr;
elsif nramp = '0' and StoredData = "110100010101" then SHout <= '1' after delay1 + 3349*delay_incr;
elsif nramp = '0' and StoredData = "110100010110" then SHout <= '1' after delay1 + 3350*delay_incr;
elsif nramp = '0' and StoredData = "110100010111" then SHout <= '1' after delay1 + 3351*delay_incr;
elsif nramp = '0' and StoredData = "110100011000" then SHout <= '1' after delay1 + 3352*delay_incr;
elsif nramp = '0' and StoredData = "110100011001" then SHout <= '1' after delay1 + 3353*delay_incr;
elsif nramp = '0' and StoredData = "110100011010" then SHout <= '1' after delay1 + 3354*delay_incr;
elsif nramp = '0' and StoredData = "110100011011" then SHout <= '1' after delay1 + 3355*delay_incr;
elsif nramp = '0' and StoredData = "110100011100" then SHout <= '1' after delay1 + 3356*delay_incr;
elsif nramp = '0' and StoredData = "110100011101" then SHout <= '1' after delay1 + 3357*delay_incr;
elsif nramp = '0' and StoredData = "110100011110" then SHout <= '1' after delay1 + 3358*delay_incr;
elsif nramp = '0' and StoredData = "110100011111" then SHout <= '1' after delay1 + 3359*delay_incr;
elsif nramp = '0' and StoredData = "110100100000" then SHout <= '1' after delay1 + 3360*delay_incr;
elsif nramp = '0' and StoredData = "110100100001" then SHout <= '1' after delay1 + 3361*delay_incr;
elsif nramp = '0' and StoredData = "110100100010" then SHout <= '1' after delay1 + 3362*delay_incr;
elsif nramp = '0' and StoredData = "110100100011" then SHout <= '1' after delay1 + 3363*delay_incr;
elsif nramp = '0' and StoredData = "110100100100" then SHout <= '1' after delay1 + 3364*delay_incr;
elsif nramp = '0' and StoredData = "110100100101" then SHout <= '1' after delay1 + 3365*delay_incr;
elsif nramp = '0' and StoredData = "110100100110" then SHout <= '1' after delay1 + 3366*delay_incr;
elsif nramp = '0' and StoredData = "110100100111" then SHout <= '1' after delay1 + 3367*delay_incr;
elsif nramp = '0' and StoredData = "110100101000" then SHout <= '1' after delay1 + 3368*delay_incr;
elsif nramp = '0' and StoredData = "110100101001" then SHout <= '1' after delay1 + 3369*delay_incr;
elsif nramp = '0' and StoredData = "110100101010" then SHout <= '1' after delay1 + 3370*delay_incr;
elsif nramp = '0' and StoredData = "110100101011" then SHout <= '1' after delay1 + 3371*delay_incr;
elsif nramp = '0' and StoredData = "110100101100" then SHout <= '1' after delay1 + 3372*delay_incr;
elsif nramp = '0' and StoredData = "110100101101" then SHout <= '1' after delay1 + 3373*delay_incr;
elsif nramp = '0' and StoredData = "110100101110" then SHout <= '1' after delay1 + 3374*delay_incr;
elsif nramp = '0' and StoredData = "110100101111" then SHout <= '1' after delay1 + 3375*delay_incr;
elsif nramp = '0' and StoredData = "110100110000" then SHout <= '1' after delay1 + 3376*delay_incr;
elsif nramp = '0' and StoredData = "110100110001" then SHout <= '1' after delay1 + 3377*delay_incr;
elsif nramp = '0' and StoredData = "110100110010" then SHout <= '1' after delay1 + 3378*delay_incr;
elsif nramp = '0' and StoredData = "110100110011" then SHout <= '1' after delay1 + 3379*delay_incr;
elsif nramp = '0' and StoredData = "110100110100" then SHout <= '1' after delay1 + 3380*delay_incr;
elsif nramp = '0' and StoredData = "110100110101" then SHout <= '1' after delay1 + 3381*delay_incr;
elsif nramp = '0' and StoredData = "110100110110" then SHout <= '1' after delay1 + 3382*delay_incr;
elsif nramp = '0' and StoredData = "110100110111" then SHout <= '1' after delay1 + 3383*delay_incr;
elsif nramp = '0' and StoredData = "110100111000" then SHout <= '1' after delay1 + 3384*delay_incr;
elsif nramp = '0' and StoredData = "110100111001" then SHout <= '1' after delay1 + 3385*delay_incr;
elsif nramp = '0' and StoredData = "110100111010" then SHout <= '1' after delay1 + 3386*delay_incr;
elsif nramp = '0' and StoredData = "110100111011" then SHout <= '1' after delay1 + 3387*delay_incr;
elsif nramp = '0' and StoredData = "110100111100" then SHout <= '1' after delay1 + 3388*delay_incr;
elsif nramp = '0' and StoredData = "110100111101" then SHout <= '1' after delay1 + 3389*delay_incr;
elsif nramp = '0' and StoredData = "110100111110" then SHout <= '1' after delay1 + 3390*delay_incr;
elsif nramp = '0' and StoredData = "110100111111" then SHout <= '1' after delay1 + 3391*delay_incr;
elsif nramp = '0' and StoredData = "110101000000" then SHout <= '1' after delay1 + 3392*delay_incr;
elsif nramp = '0' and StoredData = "110101000001" then SHout <= '1' after delay1 + 3393*delay_incr;
elsif nramp = '0' and StoredData = "110101000010" then SHout <= '1' after delay1 + 3394*delay_incr;
elsif nramp = '0' and StoredData = "110101000011" then SHout <= '1' after delay1 + 3395*delay_incr;
elsif nramp = '0' and StoredData = "110101000100" then SHout <= '1' after delay1 + 3396*delay_incr;
elsif nramp = '0' and StoredData = "110101000101" then SHout <= '1' after delay1 + 3397*delay_incr;
elsif nramp = '0' and StoredData = "110101000110" then SHout <= '1' after delay1 + 3398*delay_incr;
elsif nramp = '0' and StoredData = "110101000111" then SHout <= '1' after delay1 + 3399*delay_incr;
elsif nramp = '0' and StoredData = "110101001000" then SHout <= '1' after delay1 + 3400*delay_incr;
elsif nramp = '0' and StoredData = "110101001001" then SHout <= '1' after delay1 + 3401*delay_incr;
elsif nramp = '0' and StoredData = "110101001010" then SHout <= '1' after delay1 + 3402*delay_incr;
elsif nramp = '0' and StoredData = "110101001011" then SHout <= '1' after delay1 + 3403*delay_incr;
elsif nramp = '0' and StoredData = "110101001100" then SHout <= '1' after delay1 + 3404*delay_incr;
elsif nramp = '0' and StoredData = "110101001101" then SHout <= '1' after delay1 + 3405*delay_incr;
elsif nramp = '0' and StoredData = "110101001110" then SHout <= '1' after delay1 + 3406*delay_incr;
elsif nramp = '0' and StoredData = "110101001111" then SHout <= '1' after delay1 + 3407*delay_incr;
elsif nramp = '0' and StoredData = "110101010000" then SHout <= '1' after delay1 + 3408*delay_incr;
elsif nramp = '0' and StoredData = "110101010001" then SHout <= '1' after delay1 + 3409*delay_incr;
elsif nramp = '0' and StoredData = "110101010010" then SHout <= '1' after delay1 + 3410*delay_incr;
elsif nramp = '0' and StoredData = "110101010011" then SHout <= '1' after delay1 + 3411*delay_incr;
elsif nramp = '0' and StoredData = "110101010100" then SHout <= '1' after delay1 + 3412*delay_incr;
elsif nramp = '0' and StoredData = "110101010101" then SHout <= '1' after delay1 + 3413*delay_incr;
elsif nramp = '0' and StoredData = "110101010110" then SHout <= '1' after delay1 + 3414*delay_incr;
elsif nramp = '0' and StoredData = "110101010111" then SHout <= '1' after delay1 + 3415*delay_incr;
elsif nramp = '0' and StoredData = "110101011000" then SHout <= '1' after delay1 + 3416*delay_incr;
elsif nramp = '0' and StoredData = "110101011001" then SHout <= '1' after delay1 + 3417*delay_incr;
elsif nramp = '0' and StoredData = "110101011010" then SHout <= '1' after delay1 + 3418*delay_incr;
elsif nramp = '0' and StoredData = "110101011011" then SHout <= '1' after delay1 + 3419*delay_incr;
elsif nramp = '0' and StoredData = "110101011100" then SHout <= '1' after delay1 + 3420*delay_incr;
elsif nramp = '0' and StoredData = "110101011101" then SHout <= '1' after delay1 + 3421*delay_incr;
elsif nramp = '0' and StoredData = "110101011110" then SHout <= '1' after delay1 + 3422*delay_incr;
elsif nramp = '0' and StoredData = "110101011111" then SHout <= '1' after delay1 + 3423*delay_incr;
elsif nramp = '0' and StoredData = "110101100000" then SHout <= '1' after delay1 + 3424*delay_incr;
elsif nramp = '0' and StoredData = "110101100001" then SHout <= '1' after delay1 + 3425*delay_incr;
elsif nramp = '0' and StoredData = "110101100010" then SHout <= '1' after delay1 + 3426*delay_incr;
elsif nramp = '0' and StoredData = "110101100011" then SHout <= '1' after delay1 + 3427*delay_incr;
elsif nramp = '0' and StoredData = "110101100100" then SHout <= '1' after delay1 + 3428*delay_incr;
elsif nramp = '0' and StoredData = "110101100101" then SHout <= '1' after delay1 + 3429*delay_incr;
elsif nramp = '0' and StoredData = "110101100110" then SHout <= '1' after delay1 + 3430*delay_incr;
elsif nramp = '0' and StoredData = "110101100111" then SHout <= '1' after delay1 + 3431*delay_incr;
elsif nramp = '0' and StoredData = "110101101000" then SHout <= '1' after delay1 + 3432*delay_incr;
elsif nramp = '0' and StoredData = "110101101001" then SHout <= '1' after delay1 + 3433*delay_incr;
elsif nramp = '0' and StoredData = "110101101010" then SHout <= '1' after delay1 + 3434*delay_incr;
elsif nramp = '0' and StoredData = "110101101011" then SHout <= '1' after delay1 + 3435*delay_incr;
elsif nramp = '0' and StoredData = "110101101100" then SHout <= '1' after delay1 + 3436*delay_incr;
elsif nramp = '0' and StoredData = "110101101101" then SHout <= '1' after delay1 + 3437*delay_incr;
elsif nramp = '0' and StoredData = "110101101110" then SHout <= '1' after delay1 + 3438*delay_incr;
elsif nramp = '0' and StoredData = "110101101111" then SHout <= '1' after delay1 + 3439*delay_incr;
elsif nramp = '0' and StoredData = "110101110000" then SHout <= '1' after delay1 + 3440*delay_incr;
elsif nramp = '0' and StoredData = "110101110001" then SHout <= '1' after delay1 + 3441*delay_incr;
elsif nramp = '0' and StoredData = "110101110010" then SHout <= '1' after delay1 + 3442*delay_incr;
elsif nramp = '0' and StoredData = "110101110011" then SHout <= '1' after delay1 + 3443*delay_incr;
elsif nramp = '0' and StoredData = "110101110100" then SHout <= '1' after delay1 + 3444*delay_incr;
elsif nramp = '0' and StoredData = "110101110101" then SHout <= '1' after delay1 + 3445*delay_incr;
elsif nramp = '0' and StoredData = "110101110110" then SHout <= '1' after delay1 + 3446*delay_incr;
elsif nramp = '0' and StoredData = "110101110111" then SHout <= '1' after delay1 + 3447*delay_incr;
elsif nramp = '0' and StoredData = "110101111000" then SHout <= '1' after delay1 + 3448*delay_incr;
elsif nramp = '0' and StoredData = "110101111001" then SHout <= '1' after delay1 + 3449*delay_incr;
elsif nramp = '0' and StoredData = "110101111010" then SHout <= '1' after delay1 + 3450*delay_incr;
elsif nramp = '0' and StoredData = "110101111011" then SHout <= '1' after delay1 + 3451*delay_incr;
elsif nramp = '0' and StoredData = "110101111100" then SHout <= '1' after delay1 + 3452*delay_incr;
elsif nramp = '0' and StoredData = "110101111101" then SHout <= '1' after delay1 + 3453*delay_incr;
elsif nramp = '0' and StoredData = "110101111110" then SHout <= '1' after delay1 + 3454*delay_incr;
elsif nramp = '0' and StoredData = "110101111111" then SHout <= '1' after delay1 + 3455*delay_incr;
elsif nramp = '0' and StoredData = "110110000000" then SHout <= '1' after delay1 + 3456*delay_incr;
elsif nramp = '0' and StoredData = "110110000001" then SHout <= '1' after delay1 + 3457*delay_incr;
elsif nramp = '0' and StoredData = "110110000010" then SHout <= '1' after delay1 + 3458*delay_incr;
elsif nramp = '0' and StoredData = "110110000011" then SHout <= '1' after delay1 + 3459*delay_incr;
elsif nramp = '0' and StoredData = "110110000100" then SHout <= '1' after delay1 + 3460*delay_incr;
elsif nramp = '0' and StoredData = "110110000101" then SHout <= '1' after delay1 + 3461*delay_incr;
elsif nramp = '0' and StoredData = "110110000110" then SHout <= '1' after delay1 + 3462*delay_incr;
elsif nramp = '0' and StoredData = "110110000111" then SHout <= '1' after delay1 + 3463*delay_incr;
elsif nramp = '0' and StoredData = "110110001000" then SHout <= '1' after delay1 + 3464*delay_incr;
elsif nramp = '0' and StoredData = "110110001001" then SHout <= '1' after delay1 + 3465*delay_incr;
elsif nramp = '0' and StoredData = "110110001010" then SHout <= '1' after delay1 + 3466*delay_incr;
elsif nramp = '0' and StoredData = "110110001011" then SHout <= '1' after delay1 + 3467*delay_incr;
elsif nramp = '0' and StoredData = "110110001100" then SHout <= '1' after delay1 + 3468*delay_incr;
elsif nramp = '0' and StoredData = "110110001101" then SHout <= '1' after delay1 + 3469*delay_incr;
elsif nramp = '0' and StoredData = "110110001110" then SHout <= '1' after delay1 + 3470*delay_incr;
elsif nramp = '0' and StoredData = "110110001111" then SHout <= '1' after delay1 + 3471*delay_incr;
elsif nramp = '0' and StoredData = "110110010000" then SHout <= '1' after delay1 + 3472*delay_incr;
elsif nramp = '0' and StoredData = "110110010001" then SHout <= '1' after delay1 + 3473*delay_incr;
elsif nramp = '0' and StoredData = "110110010010" then SHout <= '1' after delay1 + 3474*delay_incr;
elsif nramp = '0' and StoredData = "110110010011" then SHout <= '1' after delay1 + 3475*delay_incr;
elsif nramp = '0' and StoredData = "110110010100" then SHout <= '1' after delay1 + 3476*delay_incr;
elsif nramp = '0' and StoredData = "110110010101" then SHout <= '1' after delay1 + 3477*delay_incr;
elsif nramp = '0' and StoredData = "110110010110" then SHout <= '1' after delay1 + 3478*delay_incr;
elsif nramp = '0' and StoredData = "110110010111" then SHout <= '1' after delay1 + 3479*delay_incr;
elsif nramp = '0' and StoredData = "110110011000" then SHout <= '1' after delay1 + 3480*delay_incr;
elsif nramp = '0' and StoredData = "110110011001" then SHout <= '1' after delay1 + 3481*delay_incr;
elsif nramp = '0' and StoredData = "110110011010" then SHout <= '1' after delay1 + 3482*delay_incr;
elsif nramp = '0' and StoredData = "110110011011" then SHout <= '1' after delay1 + 3483*delay_incr;
elsif nramp = '0' and StoredData = "110110011100" then SHout <= '1' after delay1 + 3484*delay_incr;
elsif nramp = '0' and StoredData = "110110011101" then SHout <= '1' after delay1 + 3485*delay_incr;
elsif nramp = '0' and StoredData = "110110011110" then SHout <= '1' after delay1 + 3486*delay_incr;
elsif nramp = '0' and StoredData = "110110011111" then SHout <= '1' after delay1 + 3487*delay_incr;
elsif nramp = '0' and StoredData = "110110100000" then SHout <= '1' after delay1 + 3488*delay_incr;
elsif nramp = '0' and StoredData = "110110100001" then SHout <= '1' after delay1 + 3489*delay_incr;
elsif nramp = '0' and StoredData = "110110100010" then SHout <= '1' after delay1 + 3490*delay_incr;
elsif nramp = '0' and StoredData = "110110100011" then SHout <= '1' after delay1 + 3491*delay_incr;
elsif nramp = '0' and StoredData = "110110100100" then SHout <= '1' after delay1 + 3492*delay_incr;
elsif nramp = '0' and StoredData = "110110100101" then SHout <= '1' after delay1 + 3493*delay_incr;
elsif nramp = '0' and StoredData = "110110100110" then SHout <= '1' after delay1 + 3494*delay_incr;
elsif nramp = '0' and StoredData = "110110100111" then SHout <= '1' after delay1 + 3495*delay_incr;
elsif nramp = '0' and StoredData = "110110101000" then SHout <= '1' after delay1 + 3496*delay_incr;
elsif nramp = '0' and StoredData = "110110101001" then SHout <= '1' after delay1 + 3497*delay_incr;
elsif nramp = '0' and StoredData = "110110101010" then SHout <= '1' after delay1 + 3498*delay_incr;
elsif nramp = '0' and StoredData = "110110101011" then SHout <= '1' after delay1 + 3499*delay_incr;
elsif nramp = '0' and StoredData = "110110101100" then SHout <= '1' after delay1 + 3500*delay_incr;
elsif nramp = '0' and StoredData = "110110101101" then SHout <= '1' after delay1 + 3501*delay_incr;
elsif nramp = '0' and StoredData = "110110101110" then SHout <= '1' after delay1 + 3502*delay_incr;
elsif nramp = '0' and StoredData = "110110101111" then SHout <= '1' after delay1 + 3503*delay_incr;
elsif nramp = '0' and StoredData = "110110110000" then SHout <= '1' after delay1 + 3504*delay_incr;
elsif nramp = '0' and StoredData = "110110110001" then SHout <= '1' after delay1 + 3505*delay_incr;
elsif nramp = '0' and StoredData = "110110110010" then SHout <= '1' after delay1 + 3506*delay_incr;
elsif nramp = '0' and StoredData = "110110110011" then SHout <= '1' after delay1 + 3507*delay_incr;
elsif nramp = '0' and StoredData = "110110110100" then SHout <= '1' after delay1 + 3508*delay_incr;
elsif nramp = '0' and StoredData = "110110110101" then SHout <= '1' after delay1 + 3509*delay_incr;
elsif nramp = '0' and StoredData = "110110110110" then SHout <= '1' after delay1 + 3510*delay_incr;
elsif nramp = '0' and StoredData = "110110110111" then SHout <= '1' after delay1 + 3511*delay_incr;
elsif nramp = '0' and StoredData = "110110111000" then SHout <= '1' after delay1 + 3512*delay_incr;
elsif nramp = '0' and StoredData = "110110111001" then SHout <= '1' after delay1 + 3513*delay_incr;
elsif nramp = '0' and StoredData = "110110111010" then SHout <= '1' after delay1 + 3514*delay_incr;
elsif nramp = '0' and StoredData = "110110111011" then SHout <= '1' after delay1 + 3515*delay_incr;
elsif nramp = '0' and StoredData = "110110111100" then SHout <= '1' after delay1 + 3516*delay_incr;
elsif nramp = '0' and StoredData = "110110111101" then SHout <= '1' after delay1 + 3517*delay_incr;
elsif nramp = '0' and StoredData = "110110111110" then SHout <= '1' after delay1 + 3518*delay_incr;
elsif nramp = '0' and StoredData = "110110111111" then SHout <= '1' after delay1 + 3519*delay_incr;
elsif nramp = '0' and StoredData = "110111000000" then SHout <= '1' after delay1 + 3520*delay_incr;
elsif nramp = '0' and StoredData = "110111000001" then SHout <= '1' after delay1 + 3521*delay_incr;
elsif nramp = '0' and StoredData = "110111000010" then SHout <= '1' after delay1 + 3522*delay_incr;
elsif nramp = '0' and StoredData = "110111000011" then SHout <= '1' after delay1 + 3523*delay_incr;
elsif nramp = '0' and StoredData = "110111000100" then SHout <= '1' after delay1 + 3524*delay_incr;
elsif nramp = '0' and StoredData = "110111000101" then SHout <= '1' after delay1 + 3525*delay_incr;
elsif nramp = '0' and StoredData = "110111000110" then SHout <= '1' after delay1 + 3526*delay_incr;
elsif nramp = '0' and StoredData = "110111000111" then SHout <= '1' after delay1 + 3527*delay_incr;
elsif nramp = '0' and StoredData = "110111001000" then SHout <= '1' after delay1 + 3528*delay_incr;
elsif nramp = '0' and StoredData = "110111001001" then SHout <= '1' after delay1 + 3529*delay_incr;
elsif nramp = '0' and StoredData = "110111001010" then SHout <= '1' after delay1 + 3530*delay_incr;
elsif nramp = '0' and StoredData = "110111001011" then SHout <= '1' after delay1 + 3531*delay_incr;
elsif nramp = '0' and StoredData = "110111001100" then SHout <= '1' after delay1 + 3532*delay_incr;
elsif nramp = '0' and StoredData = "110111001101" then SHout <= '1' after delay1 + 3533*delay_incr;
elsif nramp = '0' and StoredData = "110111001110" then SHout <= '1' after delay1 + 3534*delay_incr;
elsif nramp = '0' and StoredData = "110111001111" then SHout <= '1' after delay1 + 3535*delay_incr;
elsif nramp = '0' and StoredData = "110111010000" then SHout <= '1' after delay1 + 3536*delay_incr;
elsif nramp = '0' and StoredData = "110111010001" then SHout <= '1' after delay1 + 3537*delay_incr;
elsif nramp = '0' and StoredData = "110111010010" then SHout <= '1' after delay1 + 3538*delay_incr;
elsif nramp = '0' and StoredData = "110111010011" then SHout <= '1' after delay1 + 3539*delay_incr;
elsif nramp = '0' and StoredData = "110111010100" then SHout <= '1' after delay1 + 3540*delay_incr;
elsif nramp = '0' and StoredData = "110111010101" then SHout <= '1' after delay1 + 3541*delay_incr;
elsif nramp = '0' and StoredData = "110111010110" then SHout <= '1' after delay1 + 3542*delay_incr;
elsif nramp = '0' and StoredData = "110111010111" then SHout <= '1' after delay1 + 3543*delay_incr;
elsif nramp = '0' and StoredData = "110111011000" then SHout <= '1' after delay1 + 3544*delay_incr;
elsif nramp = '0' and StoredData = "110111011001" then SHout <= '1' after delay1 + 3545*delay_incr;
elsif nramp = '0' and StoredData = "110111011010" then SHout <= '1' after delay1 + 3546*delay_incr;
elsif nramp = '0' and StoredData = "110111011011" then SHout <= '1' after delay1 + 3547*delay_incr;
elsif nramp = '0' and StoredData = "110111011100" then SHout <= '1' after delay1 + 3548*delay_incr;
elsif nramp = '0' and StoredData = "110111011101" then SHout <= '1' after delay1 + 3549*delay_incr;
elsif nramp = '0' and StoredData = "110111011110" then SHout <= '1' after delay1 + 3550*delay_incr;
elsif nramp = '0' and StoredData = "110111011111" then SHout <= '1' after delay1 + 3551*delay_incr;
elsif nramp = '0' and StoredData = "110111100000" then SHout <= '1' after delay1 + 3552*delay_incr;
elsif nramp = '0' and StoredData = "110111100001" then SHout <= '1' after delay1 + 3553*delay_incr;
elsif nramp = '0' and StoredData = "110111100010" then SHout <= '1' after delay1 + 3554*delay_incr;
elsif nramp = '0' and StoredData = "110111100011" then SHout <= '1' after delay1 + 3555*delay_incr;
elsif nramp = '0' and StoredData = "110111100100" then SHout <= '1' after delay1 + 3556*delay_incr;
elsif nramp = '0' and StoredData = "110111100101" then SHout <= '1' after delay1 + 3557*delay_incr;
elsif nramp = '0' and StoredData = "110111100110" then SHout <= '1' after delay1 + 3558*delay_incr;
elsif nramp = '0' and StoredData = "110111100111" then SHout <= '1' after delay1 + 3559*delay_incr;
elsif nramp = '0' and StoredData = "110111101000" then SHout <= '1' after delay1 + 3560*delay_incr;
elsif nramp = '0' and StoredData = "110111101001" then SHout <= '1' after delay1 + 3561*delay_incr;
elsif nramp = '0' and StoredData = "110111101010" then SHout <= '1' after delay1 + 3562*delay_incr;
elsif nramp = '0' and StoredData = "110111101011" then SHout <= '1' after delay1 + 3563*delay_incr;
elsif nramp = '0' and StoredData = "110111101100" then SHout <= '1' after delay1 + 3564*delay_incr;
elsif nramp = '0' and StoredData = "110111101101" then SHout <= '1' after delay1 + 3565*delay_incr;
elsif nramp = '0' and StoredData = "110111101110" then SHout <= '1' after delay1 + 3566*delay_incr;
elsif nramp = '0' and StoredData = "110111101111" then SHout <= '1' after delay1 + 3567*delay_incr;
elsif nramp = '0' and StoredData = "110111110000" then SHout <= '1' after delay1 + 3568*delay_incr;
elsif nramp = '0' and StoredData = "110111110001" then SHout <= '1' after delay1 + 3569*delay_incr;
elsif nramp = '0' and StoredData = "110111110010" then SHout <= '1' after delay1 + 3570*delay_incr;
elsif nramp = '0' and StoredData = "110111110011" then SHout <= '1' after delay1 + 3571*delay_incr;
elsif nramp = '0' and StoredData = "110111110100" then SHout <= '1' after delay1 + 3572*delay_incr;
elsif nramp = '0' and StoredData = "110111110101" then SHout <= '1' after delay1 + 3573*delay_incr;
elsif nramp = '0' and StoredData = "110111110110" then SHout <= '1' after delay1 + 3574*delay_incr;
elsif nramp = '0' and StoredData = "110111110111" then SHout <= '1' after delay1 + 3575*delay_incr;
elsif nramp = '0' and StoredData = "110111111000" then SHout <= '1' after delay1 + 3576*delay_incr;
elsif nramp = '0' and StoredData = "110111111001" then SHout <= '1' after delay1 + 3577*delay_incr;
elsif nramp = '0' and StoredData = "110111111010" then SHout <= '1' after delay1 + 3578*delay_incr;
elsif nramp = '0' and StoredData = "110111111011" then SHout <= '1' after delay1 + 3579*delay_incr;
elsif nramp = '0' and StoredData = "110111111100" then SHout <= '1' after delay1 + 3580*delay_incr;
elsif nramp = '0' and StoredData = "110111111101" then SHout <= '1' after delay1 + 3581*delay_incr;
elsif nramp = '0' and StoredData = "110111111110" then SHout <= '1' after delay1 + 3582*delay_incr;
elsif nramp = '0' and StoredData = "110111111111" then SHout <= '1' after delay1 + 3583*delay_incr;
elsif nramp = '0' and StoredData = "111000000000" then SHout <= '1' after delay1 + 3584*delay_incr;
elsif nramp = '0' and StoredData = "111000000001" then SHout <= '1' after delay1 + 3585*delay_incr;
elsif nramp = '0' and StoredData = "111000000010" then SHout <= '1' after delay1 + 3586*delay_incr;
elsif nramp = '0' and StoredData = "111000000011" then SHout <= '1' after delay1 + 3587*delay_incr;
elsif nramp = '0' and StoredData = "111000000100" then SHout <= '1' after delay1 + 3588*delay_incr;
elsif nramp = '0' and StoredData = "111000000101" then SHout <= '1' after delay1 + 3589*delay_incr;
elsif nramp = '0' and StoredData = "111000000110" then SHout <= '1' after delay1 + 3590*delay_incr;
elsif nramp = '0' and StoredData = "111000000111" then SHout <= '1' after delay1 + 3591*delay_incr;
elsif nramp = '0' and StoredData = "111000001000" then SHout <= '1' after delay1 + 3592*delay_incr;
elsif nramp = '0' and StoredData = "111000001001" then SHout <= '1' after delay1 + 3593*delay_incr;
elsif nramp = '0' and StoredData = "111000001010" then SHout <= '1' after delay1 + 3594*delay_incr;
elsif nramp = '0' and StoredData = "111000001011" then SHout <= '1' after delay1 + 3595*delay_incr;
elsif nramp = '0' and StoredData = "111000001100" then SHout <= '1' after delay1 + 3596*delay_incr;
elsif nramp = '0' and StoredData = "111000001101" then SHout <= '1' after delay1 + 3597*delay_incr;
elsif nramp = '0' and StoredData = "111000001110" then SHout <= '1' after delay1 + 3598*delay_incr;
elsif nramp = '0' and StoredData = "111000001111" then SHout <= '1' after delay1 + 3599*delay_incr;
elsif nramp = '0' and StoredData = "111000010000" then SHout <= '1' after delay1 + 3600*delay_incr;
elsif nramp = '0' and StoredData = "111000010001" then SHout <= '1' after delay1 + 3601*delay_incr;
elsif nramp = '0' and StoredData = "111000010010" then SHout <= '1' after delay1 + 3602*delay_incr;
elsif nramp = '0' and StoredData = "111000010011" then SHout <= '1' after delay1 + 3603*delay_incr;
elsif nramp = '0' and StoredData = "111000010100" then SHout <= '1' after delay1 + 3604*delay_incr;
elsif nramp = '0' and StoredData = "111000010101" then SHout <= '1' after delay1 + 3605*delay_incr;
elsif nramp = '0' and StoredData = "111000010110" then SHout <= '1' after delay1 + 3606*delay_incr;
elsif nramp = '0' and StoredData = "111000010111" then SHout <= '1' after delay1 + 3607*delay_incr;
elsif nramp = '0' and StoredData = "111000011000" then SHout <= '1' after delay1 + 3608*delay_incr;
elsif nramp = '0' and StoredData = "111000011001" then SHout <= '1' after delay1 + 3609*delay_incr;
elsif nramp = '0' and StoredData = "111000011010" then SHout <= '1' after delay1 + 3610*delay_incr;
elsif nramp = '0' and StoredData = "111000011011" then SHout <= '1' after delay1 + 3611*delay_incr;
elsif nramp = '0' and StoredData = "111000011100" then SHout <= '1' after delay1 + 3612*delay_incr;
elsif nramp = '0' and StoredData = "111000011101" then SHout <= '1' after delay1 + 3613*delay_incr;
elsif nramp = '0' and StoredData = "111000011110" then SHout <= '1' after delay1 + 3614*delay_incr;
elsif nramp = '0' and StoredData = "111000011111" then SHout <= '1' after delay1 + 3615*delay_incr;
elsif nramp = '0' and StoredData = "111000100000" then SHout <= '1' after delay1 + 3616*delay_incr;
elsif nramp = '0' and StoredData = "111000100001" then SHout <= '1' after delay1 + 3617*delay_incr;
elsif nramp = '0' and StoredData = "111000100010" then SHout <= '1' after delay1 + 3618*delay_incr;
elsif nramp = '0' and StoredData = "111000100011" then SHout <= '1' after delay1 + 3619*delay_incr;
elsif nramp = '0' and StoredData = "111000100100" then SHout <= '1' after delay1 + 3620*delay_incr;
elsif nramp = '0' and StoredData = "111000100101" then SHout <= '1' after delay1 + 3621*delay_incr;
elsif nramp = '0' and StoredData = "111000100110" then SHout <= '1' after delay1 + 3622*delay_incr;
elsif nramp = '0' and StoredData = "111000100111" then SHout <= '1' after delay1 + 3623*delay_incr;
elsif nramp = '0' and StoredData = "111000101000" then SHout <= '1' after delay1 + 3624*delay_incr;
elsif nramp = '0' and StoredData = "111000101001" then SHout <= '1' after delay1 + 3625*delay_incr;
elsif nramp = '0' and StoredData = "111000101010" then SHout <= '1' after delay1 + 3626*delay_incr;
elsif nramp = '0' and StoredData = "111000101011" then SHout <= '1' after delay1 + 3627*delay_incr;
elsif nramp = '0' and StoredData = "111000101100" then SHout <= '1' after delay1 + 3628*delay_incr;
elsif nramp = '0' and StoredData = "111000101101" then SHout <= '1' after delay1 + 3629*delay_incr;
elsif nramp = '0' and StoredData = "111000101110" then SHout <= '1' after delay1 + 3630*delay_incr;
elsif nramp = '0' and StoredData = "111000101111" then SHout <= '1' after delay1 + 3631*delay_incr;
elsif nramp = '0' and StoredData = "111000110000" then SHout <= '1' after delay1 + 3632*delay_incr;
elsif nramp = '0' and StoredData = "111000110001" then SHout <= '1' after delay1 + 3633*delay_incr;
elsif nramp = '0' and StoredData = "111000110010" then SHout <= '1' after delay1 + 3634*delay_incr;
elsif nramp = '0' and StoredData = "111000110011" then SHout <= '1' after delay1 + 3635*delay_incr;
elsif nramp = '0' and StoredData = "111000110100" then SHout <= '1' after delay1 + 3636*delay_incr;
elsif nramp = '0' and StoredData = "111000110101" then SHout <= '1' after delay1 + 3637*delay_incr;
elsif nramp = '0' and StoredData = "111000110110" then SHout <= '1' after delay1 + 3638*delay_incr;
elsif nramp = '0' and StoredData = "111000110111" then SHout <= '1' after delay1 + 3639*delay_incr;
elsif nramp = '0' and StoredData = "111000111000" then SHout <= '1' after delay1 + 3640*delay_incr;
elsif nramp = '0' and StoredData = "111000111001" then SHout <= '1' after delay1 + 3641*delay_incr;
elsif nramp = '0' and StoredData = "111000111010" then SHout <= '1' after delay1 + 3642*delay_incr;
elsif nramp = '0' and StoredData = "111000111011" then SHout <= '1' after delay1 + 3643*delay_incr;
elsif nramp = '0' and StoredData = "111000111100" then SHout <= '1' after delay1 + 3644*delay_incr;
elsif nramp = '0' and StoredData = "111000111101" then SHout <= '1' after delay1 + 3645*delay_incr;
elsif nramp = '0' and StoredData = "111000111110" then SHout <= '1' after delay1 + 3646*delay_incr;
elsif nramp = '0' and StoredData = "111000111111" then SHout <= '1' after delay1 + 3647*delay_incr;
elsif nramp = '0' and StoredData = "111001000000" then SHout <= '1' after delay1 + 3648*delay_incr;
elsif nramp = '0' and StoredData = "111001000001" then SHout <= '1' after delay1 + 3649*delay_incr;
elsif nramp = '0' and StoredData = "111001000010" then SHout <= '1' after delay1 + 3650*delay_incr;
elsif nramp = '0' and StoredData = "111001000011" then SHout <= '1' after delay1 + 3651*delay_incr;
elsif nramp = '0' and StoredData = "111001000100" then SHout <= '1' after delay1 + 3652*delay_incr;
elsif nramp = '0' and StoredData = "111001000101" then SHout <= '1' after delay1 + 3653*delay_incr;
elsif nramp = '0' and StoredData = "111001000110" then SHout <= '1' after delay1 + 3654*delay_incr;
elsif nramp = '0' and StoredData = "111001000111" then SHout <= '1' after delay1 + 3655*delay_incr;
elsif nramp = '0' and StoredData = "111001001000" then SHout <= '1' after delay1 + 3656*delay_incr;
elsif nramp = '0' and StoredData = "111001001001" then SHout <= '1' after delay1 + 3657*delay_incr;
elsif nramp = '0' and StoredData = "111001001010" then SHout <= '1' after delay1 + 3658*delay_incr;
elsif nramp = '0' and StoredData = "111001001011" then SHout <= '1' after delay1 + 3659*delay_incr;
elsif nramp = '0' and StoredData = "111001001100" then SHout <= '1' after delay1 + 3660*delay_incr;
elsif nramp = '0' and StoredData = "111001001101" then SHout <= '1' after delay1 + 3661*delay_incr;
elsif nramp = '0' and StoredData = "111001001110" then SHout <= '1' after delay1 + 3662*delay_incr;
elsif nramp = '0' and StoredData = "111001001111" then SHout <= '1' after delay1 + 3663*delay_incr;
elsif nramp = '0' and StoredData = "111001010000" then SHout <= '1' after delay1 + 3664*delay_incr;
elsif nramp = '0' and StoredData = "111001010001" then SHout <= '1' after delay1 + 3665*delay_incr;
elsif nramp = '0' and StoredData = "111001010010" then SHout <= '1' after delay1 + 3666*delay_incr;
elsif nramp = '0' and StoredData = "111001010011" then SHout <= '1' after delay1 + 3667*delay_incr;
elsif nramp = '0' and StoredData = "111001010100" then SHout <= '1' after delay1 + 3668*delay_incr;
elsif nramp = '0' and StoredData = "111001010101" then SHout <= '1' after delay1 + 3669*delay_incr;
elsif nramp = '0' and StoredData = "111001010110" then SHout <= '1' after delay1 + 3670*delay_incr;
elsif nramp = '0' and StoredData = "111001010111" then SHout <= '1' after delay1 + 3671*delay_incr;
elsif nramp = '0' and StoredData = "111001011000" then SHout <= '1' after delay1 + 3672*delay_incr;
elsif nramp = '0' and StoredData = "111001011001" then SHout <= '1' after delay1 + 3673*delay_incr;
elsif nramp = '0' and StoredData = "111001011010" then SHout <= '1' after delay1 + 3674*delay_incr;
elsif nramp = '0' and StoredData = "111001011011" then SHout <= '1' after delay1 + 3675*delay_incr;
elsif nramp = '0' and StoredData = "111001011100" then SHout <= '1' after delay1 + 3676*delay_incr;
elsif nramp = '0' and StoredData = "111001011101" then SHout <= '1' after delay1 + 3677*delay_incr;
elsif nramp = '0' and StoredData = "111001011110" then SHout <= '1' after delay1 + 3678*delay_incr;
elsif nramp = '0' and StoredData = "111001011111" then SHout <= '1' after delay1 + 3679*delay_incr;
elsif nramp = '0' and StoredData = "111001100000" then SHout <= '1' after delay1 + 3680*delay_incr;
elsif nramp = '0' and StoredData = "111001100001" then SHout <= '1' after delay1 + 3681*delay_incr;
elsif nramp = '0' and StoredData = "111001100010" then SHout <= '1' after delay1 + 3682*delay_incr;
elsif nramp = '0' and StoredData = "111001100011" then SHout <= '1' after delay1 + 3683*delay_incr;
elsif nramp = '0' and StoredData = "111001100100" then SHout <= '1' after delay1 + 3684*delay_incr;
elsif nramp = '0' and StoredData = "111001100101" then SHout <= '1' after delay1 + 3685*delay_incr;
elsif nramp = '0' and StoredData = "111001100110" then SHout <= '1' after delay1 + 3686*delay_incr;
elsif nramp = '0' and StoredData = "111001100111" then SHout <= '1' after delay1 + 3687*delay_incr;
elsif nramp = '0' and StoredData = "111001101000" then SHout <= '1' after delay1 + 3688*delay_incr;
elsif nramp = '0' and StoredData = "111001101001" then SHout <= '1' after delay1 + 3689*delay_incr;
elsif nramp = '0' and StoredData = "111001101010" then SHout <= '1' after delay1 + 3690*delay_incr;
elsif nramp = '0' and StoredData = "111001101011" then SHout <= '1' after delay1 + 3691*delay_incr;
elsif nramp = '0' and StoredData = "111001101100" then SHout <= '1' after delay1 + 3692*delay_incr;
elsif nramp = '0' and StoredData = "111001101101" then SHout <= '1' after delay1 + 3693*delay_incr;
elsif nramp = '0' and StoredData = "111001101110" then SHout <= '1' after delay1 + 3694*delay_incr;
elsif nramp = '0' and StoredData = "111001101111" then SHout <= '1' after delay1 + 3695*delay_incr;
elsif nramp = '0' and StoredData = "111001110000" then SHout <= '1' after delay1 + 3696*delay_incr;
elsif nramp = '0' and StoredData = "111001110001" then SHout <= '1' after delay1 + 3697*delay_incr;
elsif nramp = '0' and StoredData = "111001110010" then SHout <= '1' after delay1 + 3698*delay_incr;
elsif nramp = '0' and StoredData = "111001110011" then SHout <= '1' after delay1 + 3699*delay_incr;
elsif nramp = '0' and StoredData = "111001110100" then SHout <= '1' after delay1 + 3700*delay_incr;
elsif nramp = '0' and StoredData = "111001110101" then SHout <= '1' after delay1 + 3701*delay_incr;
elsif nramp = '0' and StoredData = "111001110110" then SHout <= '1' after delay1 + 3702*delay_incr;
elsif nramp = '0' and StoredData = "111001110111" then SHout <= '1' after delay1 + 3703*delay_incr;
elsif nramp = '0' and StoredData = "111001111000" then SHout <= '1' after delay1 + 3704*delay_incr;
elsif nramp = '0' and StoredData = "111001111001" then SHout <= '1' after delay1 + 3705*delay_incr;
elsif nramp = '0' and StoredData = "111001111010" then SHout <= '1' after delay1 + 3706*delay_incr;
elsif nramp = '0' and StoredData = "111001111011" then SHout <= '1' after delay1 + 3707*delay_incr;
elsif nramp = '0' and StoredData = "111001111100" then SHout <= '1' after delay1 + 3708*delay_incr;
elsif nramp = '0' and StoredData = "111001111101" then SHout <= '1' after delay1 + 3709*delay_incr;
elsif nramp = '0' and StoredData = "111001111110" then SHout <= '1' after delay1 + 3710*delay_incr;
elsif nramp = '0' and StoredData = "111001111111" then SHout <= '1' after delay1 + 3711*delay_incr;
elsif nramp = '0' and StoredData = "111010000000" then SHout <= '1' after delay1 + 3712*delay_incr;
elsif nramp = '0' and StoredData = "111010000001" then SHout <= '1' after delay1 + 3713*delay_incr;
elsif nramp = '0' and StoredData = "111010000010" then SHout <= '1' after delay1 + 3714*delay_incr;
elsif nramp = '0' and StoredData = "111010000011" then SHout <= '1' after delay1 + 3715*delay_incr;
elsif nramp = '0' and StoredData = "111010000100" then SHout <= '1' after delay1 + 3716*delay_incr;
elsif nramp = '0' and StoredData = "111010000101" then SHout <= '1' after delay1 + 3717*delay_incr;
elsif nramp = '0' and StoredData = "111010000110" then SHout <= '1' after delay1 + 3718*delay_incr;
elsif nramp = '0' and StoredData = "111010000111" then SHout <= '1' after delay1 + 3719*delay_incr;
elsif nramp = '0' and StoredData = "111010001000" then SHout <= '1' after delay1 + 3720*delay_incr;
elsif nramp = '0' and StoredData = "111010001001" then SHout <= '1' after delay1 + 3721*delay_incr;
elsif nramp = '0' and StoredData = "111010001010" then SHout <= '1' after delay1 + 3722*delay_incr;
elsif nramp = '0' and StoredData = "111010001011" then SHout <= '1' after delay1 + 3723*delay_incr;
elsif nramp = '0' and StoredData = "111010001100" then SHout <= '1' after delay1 + 3724*delay_incr;
elsif nramp = '0' and StoredData = "111010001101" then SHout <= '1' after delay1 + 3725*delay_incr;
elsif nramp = '0' and StoredData = "111010001110" then SHout <= '1' after delay1 + 3726*delay_incr;
elsif nramp = '0' and StoredData = "111010001111" then SHout <= '1' after delay1 + 3727*delay_incr;
elsif nramp = '0' and StoredData = "111010010000" then SHout <= '1' after delay1 + 3728*delay_incr;
elsif nramp = '0' and StoredData = "111010010001" then SHout <= '1' after delay1 + 3729*delay_incr;
elsif nramp = '0' and StoredData = "111010010010" then SHout <= '1' after delay1 + 3730*delay_incr;
elsif nramp = '0' and StoredData = "111010010011" then SHout <= '1' after delay1 + 3731*delay_incr;
elsif nramp = '0' and StoredData = "111010010100" then SHout <= '1' after delay1 + 3732*delay_incr;
elsif nramp = '0' and StoredData = "111010010101" then SHout <= '1' after delay1 + 3733*delay_incr;
elsif nramp = '0' and StoredData = "111010010110" then SHout <= '1' after delay1 + 3734*delay_incr;
elsif nramp = '0' and StoredData = "111010010111" then SHout <= '1' after delay1 + 3735*delay_incr;
elsif nramp = '0' and StoredData = "111010011000" then SHout <= '1' after delay1 + 3736*delay_incr;
elsif nramp = '0' and StoredData = "111010011001" then SHout <= '1' after delay1 + 3737*delay_incr;
elsif nramp = '0' and StoredData = "111010011010" then SHout <= '1' after delay1 + 3738*delay_incr;
elsif nramp = '0' and StoredData = "111010011011" then SHout <= '1' after delay1 + 3739*delay_incr;
elsif nramp = '0' and StoredData = "111010011100" then SHout <= '1' after delay1 + 3740*delay_incr;
elsif nramp = '0' and StoredData = "111010011101" then SHout <= '1' after delay1 + 3741*delay_incr;
elsif nramp = '0' and StoredData = "111010011110" then SHout <= '1' after delay1 + 3742*delay_incr;
elsif nramp = '0' and StoredData = "111010011111" then SHout <= '1' after delay1 + 3743*delay_incr;
elsif nramp = '0' and StoredData = "111010100000" then SHout <= '1' after delay1 + 3744*delay_incr;
elsif nramp = '0' and StoredData = "111010100001" then SHout <= '1' after delay1 + 3745*delay_incr;
elsif nramp = '0' and StoredData = "111010100010" then SHout <= '1' after delay1 + 3746*delay_incr;
elsif nramp = '0' and StoredData = "111010100011" then SHout <= '1' after delay1 + 3747*delay_incr;
elsif nramp = '0' and StoredData = "111010100100" then SHout <= '1' after delay1 + 3748*delay_incr;
elsif nramp = '0' and StoredData = "111010100101" then SHout <= '1' after delay1 + 3749*delay_incr;
elsif nramp = '0' and StoredData = "111010100110" then SHout <= '1' after delay1 + 3750*delay_incr;
elsif nramp = '0' and StoredData = "111010100111" then SHout <= '1' after delay1 + 3751*delay_incr;
elsif nramp = '0' and StoredData = "111010101000" then SHout <= '1' after delay1 + 3752*delay_incr;
elsif nramp = '0' and StoredData = "111010101001" then SHout <= '1' after delay1 + 3753*delay_incr;
elsif nramp = '0' and StoredData = "111010101010" then SHout <= '1' after delay1 + 3754*delay_incr;
elsif nramp = '0' and StoredData = "111010101011" then SHout <= '1' after delay1 + 3755*delay_incr;
elsif nramp = '0' and StoredData = "111010101100" then SHout <= '1' after delay1 + 3756*delay_incr;
elsif nramp = '0' and StoredData = "111010101101" then SHout <= '1' after delay1 + 3757*delay_incr;
elsif nramp = '0' and StoredData = "111010101110" then SHout <= '1' after delay1 + 3758*delay_incr;
elsif nramp = '0' and StoredData = "111010101111" then SHout <= '1' after delay1 + 3759*delay_incr;
elsif nramp = '0' and StoredData = "111010110000" then SHout <= '1' after delay1 + 3760*delay_incr;
elsif nramp = '0' and StoredData = "111010110001" then SHout <= '1' after delay1 + 3761*delay_incr;
elsif nramp = '0' and StoredData = "111010110010" then SHout <= '1' after delay1 + 3762*delay_incr;
elsif nramp = '0' and StoredData = "111010110011" then SHout <= '1' after delay1 + 3763*delay_incr;
elsif nramp = '0' and StoredData = "111010110100" then SHout <= '1' after delay1 + 3764*delay_incr;
elsif nramp = '0' and StoredData = "111010110101" then SHout <= '1' after delay1 + 3765*delay_incr;
elsif nramp = '0' and StoredData = "111010110110" then SHout <= '1' after delay1 + 3766*delay_incr;
elsif nramp = '0' and StoredData = "111010110111" then SHout <= '1' after delay1 + 3767*delay_incr;
elsif nramp = '0' and StoredData = "111010111000" then SHout <= '1' after delay1 + 3768*delay_incr;
elsif nramp = '0' and StoredData = "111010111001" then SHout <= '1' after delay1 + 3769*delay_incr;
elsif nramp = '0' and StoredData = "111010111010" then SHout <= '1' after delay1 + 3770*delay_incr;
elsif nramp = '0' and StoredData = "111010111011" then SHout <= '1' after delay1 + 3771*delay_incr;
elsif nramp = '0' and StoredData = "111010111100" then SHout <= '1' after delay1 + 3772*delay_incr;
elsif nramp = '0' and StoredData = "111010111101" then SHout <= '1' after delay1 + 3773*delay_incr;
elsif nramp = '0' and StoredData = "111010111110" then SHout <= '1' after delay1 + 3774*delay_incr;
elsif nramp = '0' and StoredData = "111010111111" then SHout <= '1' after delay1 + 3775*delay_incr;
elsif nramp = '0' and StoredData = "111011000000" then SHout <= '1' after delay1 + 3776*delay_incr;
elsif nramp = '0' and StoredData = "111011000001" then SHout <= '1' after delay1 + 3777*delay_incr;
elsif nramp = '0' and StoredData = "111011000010" then SHout <= '1' after delay1 + 3778*delay_incr;
elsif nramp = '0' and StoredData = "111011000011" then SHout <= '1' after delay1 + 3779*delay_incr;
elsif nramp = '0' and StoredData = "111011000100" then SHout <= '1' after delay1 + 3780*delay_incr;
elsif nramp = '0' and StoredData = "111011000101" then SHout <= '1' after delay1 + 3781*delay_incr;
elsif nramp = '0' and StoredData = "111011000110" then SHout <= '1' after delay1 + 3782*delay_incr;
elsif nramp = '0' and StoredData = "111011000111" then SHout <= '1' after delay1 + 3783*delay_incr;
elsif nramp = '0' and StoredData = "111011001000" then SHout <= '1' after delay1 + 3784*delay_incr;
elsif nramp = '0' and StoredData = "111011001001" then SHout <= '1' after delay1 + 3785*delay_incr;
elsif nramp = '0' and StoredData = "111011001010" then SHout <= '1' after delay1 + 3786*delay_incr;
elsif nramp = '0' and StoredData = "111011001011" then SHout <= '1' after delay1 + 3787*delay_incr;
elsif nramp = '0' and StoredData = "111011001100" then SHout <= '1' after delay1 + 3788*delay_incr;
elsif nramp = '0' and StoredData = "111011001101" then SHout <= '1' after delay1 + 3789*delay_incr;
elsif nramp = '0' and StoredData = "111011001110" then SHout <= '1' after delay1 + 3790*delay_incr;
elsif nramp = '0' and StoredData = "111011001111" then SHout <= '1' after delay1 + 3791*delay_incr;
elsif nramp = '0' and StoredData = "111011010000" then SHout <= '1' after delay1 + 3792*delay_incr;
elsif nramp = '0' and StoredData = "111011010001" then SHout <= '1' after delay1 + 3793*delay_incr;
elsif nramp = '0' and StoredData = "111011010010" then SHout <= '1' after delay1 + 3794*delay_incr;
elsif nramp = '0' and StoredData = "111011010011" then SHout <= '1' after delay1 + 3795*delay_incr;
elsif nramp = '0' and StoredData = "111011010100" then SHout <= '1' after delay1 + 3796*delay_incr;
elsif nramp = '0' and StoredData = "111011010101" then SHout <= '1' after delay1 + 3797*delay_incr;
elsif nramp = '0' and StoredData = "111011010110" then SHout <= '1' after delay1 + 3798*delay_incr;
elsif nramp = '0' and StoredData = "111011010111" then SHout <= '1' after delay1 + 3799*delay_incr;
elsif nramp = '0' and StoredData = "111011011000" then SHout <= '1' after delay1 + 3800*delay_incr;
elsif nramp = '0' and StoredData = "111011011001" then SHout <= '1' after delay1 + 3801*delay_incr;
elsif nramp = '0' and StoredData = "111011011010" then SHout <= '1' after delay1 + 3802*delay_incr;
elsif nramp = '0' and StoredData = "111011011011" then SHout <= '1' after delay1 + 3803*delay_incr;
elsif nramp = '0' and StoredData = "111011011100" then SHout <= '1' after delay1 + 3804*delay_incr;
elsif nramp = '0' and StoredData = "111011011101" then SHout <= '1' after delay1 + 3805*delay_incr;
elsif nramp = '0' and StoredData = "111011011110" then SHout <= '1' after delay1 + 3806*delay_incr;
elsif nramp = '0' and StoredData = "111011011111" then SHout <= '1' after delay1 + 3807*delay_incr;
elsif nramp = '0' and StoredData = "111011100000" then SHout <= '1' after delay1 + 3808*delay_incr;
elsif nramp = '0' and StoredData = "111011100001" then SHout <= '1' after delay1 + 3809*delay_incr;
elsif nramp = '0' and StoredData = "111011100010" then SHout <= '1' after delay1 + 3810*delay_incr;
elsif nramp = '0' and StoredData = "111011100011" then SHout <= '1' after delay1 + 3811*delay_incr;
elsif nramp = '0' and StoredData = "111011100100" then SHout <= '1' after delay1 + 3812*delay_incr;
elsif nramp = '0' and StoredData = "111011100101" then SHout <= '1' after delay1 + 3813*delay_incr;
elsif nramp = '0' and StoredData = "111011100110" then SHout <= '1' after delay1 + 3814*delay_incr;
elsif nramp = '0' and StoredData = "111011100111" then SHout <= '1' after delay1 + 3815*delay_incr;
elsif nramp = '0' and StoredData = "111011101000" then SHout <= '1' after delay1 + 3816*delay_incr;
elsif nramp = '0' and StoredData = "111011101001" then SHout <= '1' after delay1 + 3817*delay_incr;
elsif nramp = '0' and StoredData = "111011101010" then SHout <= '1' after delay1 + 3818*delay_incr;
elsif nramp = '0' and StoredData = "111011101011" then SHout <= '1' after delay1 + 3819*delay_incr;
elsif nramp = '0' and StoredData = "111011101100" then SHout <= '1' after delay1 + 3820*delay_incr;
elsif nramp = '0' and StoredData = "111011101101" then SHout <= '1' after delay1 + 3821*delay_incr;
elsif nramp = '0' and StoredData = "111011101110" then SHout <= '1' after delay1 + 3822*delay_incr;
elsif nramp = '0' and StoredData = "111011101111" then SHout <= '1' after delay1 + 3823*delay_incr;
elsif nramp = '0' and StoredData = "111011110000" then SHout <= '1' after delay1 + 3824*delay_incr;
elsif nramp = '0' and StoredData = "111011110001" then SHout <= '1' after delay1 + 3825*delay_incr;
elsif nramp = '0' and StoredData = "111011110010" then SHout <= '1' after delay1 + 3826*delay_incr;
elsif nramp = '0' and StoredData = "111011110011" then SHout <= '1' after delay1 + 3827*delay_incr;
elsif nramp = '0' and StoredData = "111011110100" then SHout <= '1' after delay1 + 3828*delay_incr;
elsif nramp = '0' and StoredData = "111011110101" then SHout <= '1' after delay1 + 3829*delay_incr;
elsif nramp = '0' and StoredData = "111011110110" then SHout <= '1' after delay1 + 3830*delay_incr;
elsif nramp = '0' and StoredData = "111011110111" then SHout <= '1' after delay1 + 3831*delay_incr;
elsif nramp = '0' and StoredData = "111011111000" then SHout <= '1' after delay1 + 3832*delay_incr;
elsif nramp = '0' and StoredData = "111011111001" then SHout <= '1' after delay1 + 3833*delay_incr;
elsif nramp = '0' and StoredData = "111011111010" then SHout <= '1' after delay1 + 3834*delay_incr;
elsif nramp = '0' and StoredData = "111011111011" then SHout <= '1' after delay1 + 3835*delay_incr;
elsif nramp = '0' and StoredData = "111011111100" then SHout <= '1' after delay1 + 3836*delay_incr;
elsif nramp = '0' and StoredData = "111011111101" then SHout <= '1' after delay1 + 3837*delay_incr;
elsif nramp = '0' and StoredData = "111011111110" then SHout <= '1' after delay1 + 3838*delay_incr;
elsif nramp = '0' and StoredData = "111011111111" then SHout <= '1' after delay1 + 3839*delay_incr;
elsif nramp = '0' and StoredData = "111100000000" then SHout <= '1' after delay1 + 3840*delay_incr;
elsif nramp = '0' and StoredData = "111100000001" then SHout <= '1' after delay1 + 3841*delay_incr;
elsif nramp = '0' and StoredData = "111100000010" then SHout <= '1' after delay1 + 3842*delay_incr;
elsif nramp = '0' and StoredData = "111100000011" then SHout <= '1' after delay1 + 3843*delay_incr;
elsif nramp = '0' and StoredData = "111100000100" then SHout <= '1' after delay1 + 3844*delay_incr;
elsif nramp = '0' and StoredData = "111100000101" then SHout <= '1' after delay1 + 3845*delay_incr;
elsif nramp = '0' and StoredData = "111100000110" then SHout <= '1' after delay1 + 3846*delay_incr;
elsif nramp = '0' and StoredData = "111100000111" then SHout <= '1' after delay1 + 3847*delay_incr;
elsif nramp = '0' and StoredData = "111100001000" then SHout <= '1' after delay1 + 3848*delay_incr;
elsif nramp = '0' and StoredData = "111100001001" then SHout <= '1' after delay1 + 3849*delay_incr;
elsif nramp = '0' and StoredData = "111100001010" then SHout <= '1' after delay1 + 3850*delay_incr;
elsif nramp = '0' and StoredData = "111100001011" then SHout <= '1' after delay1 + 3851*delay_incr;
elsif nramp = '0' and StoredData = "111100001100" then SHout <= '1' after delay1 + 3852*delay_incr;
elsif nramp = '0' and StoredData = "111100001101" then SHout <= '1' after delay1 + 3853*delay_incr;
elsif nramp = '0' and StoredData = "111100001110" then SHout <= '1' after delay1 + 3854*delay_incr;
elsif nramp = '0' and StoredData = "111100001111" then SHout <= '1' after delay1 + 3855*delay_incr;
elsif nramp = '0' and StoredData = "111100010000" then SHout <= '1' after delay1 + 3856*delay_incr;
elsif nramp = '0' and StoredData = "111100010001" then SHout <= '1' after delay1 + 3857*delay_incr;
elsif nramp = '0' and StoredData = "111100010010" then SHout <= '1' after delay1 + 3858*delay_incr;
elsif nramp = '0' and StoredData = "111100010011" then SHout <= '1' after delay1 + 3859*delay_incr;
elsif nramp = '0' and StoredData = "111100010100" then SHout <= '1' after delay1 + 3860*delay_incr;
elsif nramp = '0' and StoredData = "111100010101" then SHout <= '1' after delay1 + 3861*delay_incr;
elsif nramp = '0' and StoredData = "111100010110" then SHout <= '1' after delay1 + 3862*delay_incr;
elsif nramp = '0' and StoredData = "111100010111" then SHout <= '1' after delay1 + 3863*delay_incr;
elsif nramp = '0' and StoredData = "111100011000" then SHout <= '1' after delay1 + 3864*delay_incr;
elsif nramp = '0' and StoredData = "111100011001" then SHout <= '1' after delay1 + 3865*delay_incr;
elsif nramp = '0' and StoredData = "111100011010" then SHout <= '1' after delay1 + 3866*delay_incr;
elsif nramp = '0' and StoredData = "111100011011" then SHout <= '1' after delay1 + 3867*delay_incr;
elsif nramp = '0' and StoredData = "111100011100" then SHout <= '1' after delay1 + 3868*delay_incr;
elsif nramp = '0' and StoredData = "111100011101" then SHout <= '1' after delay1 + 3869*delay_incr;
elsif nramp = '0' and StoredData = "111100011110" then SHout <= '1' after delay1 + 3870*delay_incr;
elsif nramp = '0' and StoredData = "111100011111" then SHout <= '1' after delay1 + 3871*delay_incr;
elsif nramp = '0' and StoredData = "111100100000" then SHout <= '1' after delay1 + 3872*delay_incr;
elsif nramp = '0' and StoredData = "111100100001" then SHout <= '1' after delay1 + 3873*delay_incr;
elsif nramp = '0' and StoredData = "111100100010" then SHout <= '1' after delay1 + 3874*delay_incr;
elsif nramp = '0' and StoredData = "111100100011" then SHout <= '1' after delay1 + 3875*delay_incr;
elsif nramp = '0' and StoredData = "111100100100" then SHout <= '1' after delay1 + 3876*delay_incr;
elsif nramp = '0' and StoredData = "111100100101" then SHout <= '1' after delay1 + 3877*delay_incr;
elsif nramp = '0' and StoredData = "111100100110" then SHout <= '1' after delay1 + 3878*delay_incr;
elsif nramp = '0' and StoredData = "111100100111" then SHout <= '1' after delay1 + 3879*delay_incr;
elsif nramp = '0' and StoredData = "111100101000" then SHout <= '1' after delay1 + 3880*delay_incr;
elsif nramp = '0' and StoredData = "111100101001" then SHout <= '1' after delay1 + 3881*delay_incr;
elsif nramp = '0' and StoredData = "111100101010" then SHout <= '1' after delay1 + 3882*delay_incr;
elsif nramp = '0' and StoredData = "111100101011" then SHout <= '1' after delay1 + 3883*delay_incr;
elsif nramp = '0' and StoredData = "111100101100" then SHout <= '1' after delay1 + 3884*delay_incr;
elsif nramp = '0' and StoredData = "111100101101" then SHout <= '1' after delay1 + 3885*delay_incr;
elsif nramp = '0' and StoredData = "111100101110" then SHout <= '1' after delay1 + 3886*delay_incr;
elsif nramp = '0' and StoredData = "111100101111" then SHout <= '1' after delay1 + 3887*delay_incr;
elsif nramp = '0' and StoredData = "111100110000" then SHout <= '1' after delay1 + 3888*delay_incr;
elsif nramp = '0' and StoredData = "111100110001" then SHout <= '1' after delay1 + 3889*delay_incr;
elsif nramp = '0' and StoredData = "111100110010" then SHout <= '1' after delay1 + 3890*delay_incr;
elsif nramp = '0' and StoredData = "111100110011" then SHout <= '1' after delay1 + 3891*delay_incr;
elsif nramp = '0' and StoredData = "111100110100" then SHout <= '1' after delay1 + 3892*delay_incr;
elsif nramp = '0' and StoredData = "111100110101" then SHout <= '1' after delay1 + 3893*delay_incr;
elsif nramp = '0' and StoredData = "111100110110" then SHout <= '1' after delay1 + 3894*delay_incr;
elsif nramp = '0' and StoredData = "111100110111" then SHout <= '1' after delay1 + 3895*delay_incr;
elsif nramp = '0' and StoredData = "111100111000" then SHout <= '1' after delay1 + 3896*delay_incr;
elsif nramp = '0' and StoredData = "111100111001" then SHout <= '1' after delay1 + 3897*delay_incr;
elsif nramp = '0' and StoredData = "111100111010" then SHout <= '1' after delay1 + 3898*delay_incr;
elsif nramp = '0' and StoredData = "111100111011" then SHout <= '1' after delay1 + 3899*delay_incr;
elsif nramp = '0' and StoredData = "111100111100" then SHout <= '1' after delay1 + 3900*delay_incr;
elsif nramp = '0' and StoredData = "111100111101" then SHout <= '1' after delay1 + 3901*delay_incr;
elsif nramp = '0' and StoredData = "111100111110" then SHout <= '1' after delay1 + 3902*delay_incr;
elsif nramp = '0' and StoredData = "111100111111" then SHout <= '1' after delay1 + 3903*delay_incr;
elsif nramp = '0' and StoredData = "111101000000" then SHout <= '1' after delay1 + 3904*delay_incr;
elsif nramp = '0' and StoredData = "111101000001" then SHout <= '1' after delay1 + 3905*delay_incr;
elsif nramp = '0' and StoredData = "111101000010" then SHout <= '1' after delay1 + 3906*delay_incr;
elsif nramp = '0' and StoredData = "111101000011" then SHout <= '1' after delay1 + 3907*delay_incr;
elsif nramp = '0' and StoredData = "111101000100" then SHout <= '1' after delay1 + 3908*delay_incr;
elsif nramp = '0' and StoredData = "111101000101" then SHout <= '1' after delay1 + 3909*delay_incr;
elsif nramp = '0' and StoredData = "111101000110" then SHout <= '1' after delay1 + 3910*delay_incr;
elsif nramp = '0' and StoredData = "111101000111" then SHout <= '1' after delay1 + 3911*delay_incr;
elsif nramp = '0' and StoredData = "111101001000" then SHout <= '1' after delay1 + 3912*delay_incr;
elsif nramp = '0' and StoredData = "111101001001" then SHout <= '1' after delay1 + 3913*delay_incr;
elsif nramp = '0' and StoredData = "111101001010" then SHout <= '1' after delay1 + 3914*delay_incr;
elsif nramp = '0' and StoredData = "111101001011" then SHout <= '1' after delay1 + 3915*delay_incr;
elsif nramp = '0' and StoredData = "111101001100" then SHout <= '1' after delay1 + 3916*delay_incr;
elsif nramp = '0' and StoredData = "111101001101" then SHout <= '1' after delay1 + 3917*delay_incr;
elsif nramp = '0' and StoredData = "111101001110" then SHout <= '1' after delay1 + 3918*delay_incr;
elsif nramp = '0' and StoredData = "111101001111" then SHout <= '1' after delay1 + 3919*delay_incr;
elsif nramp = '0' and StoredData = "111101010000" then SHout <= '1' after delay1 + 3920*delay_incr;
elsif nramp = '0' and StoredData = "111101010001" then SHout <= '1' after delay1 + 3921*delay_incr;
elsif nramp = '0' and StoredData = "111101010010" then SHout <= '1' after delay1 + 3922*delay_incr;
elsif nramp = '0' and StoredData = "111101010011" then SHout <= '1' after delay1 + 3923*delay_incr;
elsif nramp = '0' and StoredData = "111101010100" then SHout <= '1' after delay1 + 3924*delay_incr;
elsif nramp = '0' and StoredData = "111101010101" then SHout <= '1' after delay1 + 3925*delay_incr;
elsif nramp = '0' and StoredData = "111101010110" then SHout <= '1' after delay1 + 3926*delay_incr;
elsif nramp = '0' and StoredData = "111101010111" then SHout <= '1' after delay1 + 3927*delay_incr;
elsif nramp = '0' and StoredData = "111101011000" then SHout <= '1' after delay1 + 3928*delay_incr;
elsif nramp = '0' and StoredData = "111101011001" then SHout <= '1' after delay1 + 3929*delay_incr;
elsif nramp = '0' and StoredData = "111101011010" then SHout <= '1' after delay1 + 3930*delay_incr;
elsif nramp = '0' and StoredData = "111101011011" then SHout <= '1' after delay1 + 3931*delay_incr;
elsif nramp = '0' and StoredData = "111101011100" then SHout <= '1' after delay1 + 3932*delay_incr;
elsif nramp = '0' and StoredData = "111101011101" then SHout <= '1' after delay1 + 3933*delay_incr;
elsif nramp = '0' and StoredData = "111101011110" then SHout <= '1' after delay1 + 3934*delay_incr;
elsif nramp = '0' and StoredData = "111101011111" then SHout <= '1' after delay1 + 3935*delay_incr;
elsif nramp = '0' and StoredData = "111101100000" then SHout <= '1' after delay1 + 3936*delay_incr;
elsif nramp = '0' and StoredData = "111101100001" then SHout <= '1' after delay1 + 3937*delay_incr;
elsif nramp = '0' and StoredData = "111101100010" then SHout <= '1' after delay1 + 3938*delay_incr;
elsif nramp = '0' and StoredData = "111101100011" then SHout <= '1' after delay1 + 3939*delay_incr;
elsif nramp = '0' and StoredData = "111101100100" then SHout <= '1' after delay1 + 3940*delay_incr;
elsif nramp = '0' and StoredData = "111101100101" then SHout <= '1' after delay1 + 3941*delay_incr;
elsif nramp = '0' and StoredData = "111101100110" then SHout <= '1' after delay1 + 3942*delay_incr;
elsif nramp = '0' and StoredData = "111101100111" then SHout <= '1' after delay1 + 3943*delay_incr;
elsif nramp = '0' and StoredData = "111101101000" then SHout <= '1' after delay1 + 3944*delay_incr;
elsif nramp = '0' and StoredData = "111101101001" then SHout <= '1' after delay1 + 3945*delay_incr;
elsif nramp = '0' and StoredData = "111101101010" then SHout <= '1' after delay1 + 3946*delay_incr;
elsif nramp = '0' and StoredData = "111101101011" then SHout <= '1' after delay1 + 3947*delay_incr;
elsif nramp = '0' and StoredData = "111101101100" then SHout <= '1' after delay1 + 3948*delay_incr;
elsif nramp = '0' and StoredData = "111101101101" then SHout <= '1' after delay1 + 3949*delay_incr;
elsif nramp = '0' and StoredData = "111101101110" then SHout <= '1' after delay1 + 3950*delay_incr;
elsif nramp = '0' and StoredData = "111101101111" then SHout <= '1' after delay1 + 3951*delay_incr;
elsif nramp = '0' and StoredData = "111101110000" then SHout <= '1' after delay1 + 3952*delay_incr;
elsif nramp = '0' and StoredData = "111101110001" then SHout <= '1' after delay1 + 3953*delay_incr;
elsif nramp = '0' and StoredData = "111101110010" then SHout <= '1' after delay1 + 3954*delay_incr;
elsif nramp = '0' and StoredData = "111101110011" then SHout <= '1' after delay1 + 3955*delay_incr;
elsif nramp = '0' and StoredData = "111101110100" then SHout <= '1' after delay1 + 3956*delay_incr;
elsif nramp = '0' and StoredData = "111101110101" then SHout <= '1' after delay1 + 3957*delay_incr;
elsif nramp = '0' and StoredData = "111101110110" then SHout <= '1' after delay1 + 3958*delay_incr;
elsif nramp = '0' and StoredData = "111101110111" then SHout <= '1' after delay1 + 3959*delay_incr;
elsif nramp = '0' and StoredData = "111101111000" then SHout <= '1' after delay1 + 3960*delay_incr;
elsif nramp = '0' and StoredData = "111101111001" then SHout <= '1' after delay1 + 3961*delay_incr;
elsif nramp = '0' and StoredData = "111101111010" then SHout <= '1' after delay1 + 3962*delay_incr;
elsif nramp = '0' and StoredData = "111101111011" then SHout <= '1' after delay1 + 3963*delay_incr;
elsif nramp = '0' and StoredData = "111101111100" then SHout <= '1' after delay1 + 3964*delay_incr;
elsif nramp = '0' and StoredData = "111101111101" then SHout <= '1' after delay1 + 3965*delay_incr;
elsif nramp = '0' and StoredData = "111101111110" then SHout <= '1' after delay1 + 3966*delay_incr;
elsif nramp = '0' and StoredData = "111101111111" then SHout <= '1' after delay1 + 3967*delay_incr;
elsif nramp = '0' and StoredData = "111110000000" then SHout <= '1' after delay1 + 3968*delay_incr;
elsif nramp = '0' and StoredData = "111110000001" then SHout <= '1' after delay1 + 3969*delay_incr;
elsif nramp = '0' and StoredData = "111110000010" then SHout <= '1' after delay1 + 3970*delay_incr;
elsif nramp = '0' and StoredData = "111110000011" then SHout <= '1' after delay1 + 3971*delay_incr;
elsif nramp = '0' and StoredData = "111110000100" then SHout <= '1' after delay1 + 3972*delay_incr;
elsif nramp = '0' and StoredData = "111110000101" then SHout <= '1' after delay1 + 3973*delay_incr;
elsif nramp = '0' and StoredData = "111110000110" then SHout <= '1' after delay1 + 3974*delay_incr;
elsif nramp = '0' and StoredData = "111110000111" then SHout <= '1' after delay1 + 3975*delay_incr;
elsif nramp = '0' and StoredData = "111110001000" then SHout <= '1' after delay1 + 3976*delay_incr;
elsif nramp = '0' and StoredData = "111110001001" then SHout <= '1' after delay1 + 3977*delay_incr;
elsif nramp = '0' and StoredData = "111110001010" then SHout <= '1' after delay1 + 3978*delay_incr;
elsif nramp = '0' and StoredData = "111110001011" then SHout <= '1' after delay1 + 3979*delay_incr;
elsif nramp = '0' and StoredData = "111110001100" then SHout <= '1' after delay1 + 3980*delay_incr;
elsif nramp = '0' and StoredData = "111110001101" then SHout <= '1' after delay1 + 3981*delay_incr;
elsif nramp = '0' and StoredData = "111110001110" then SHout <= '1' after delay1 + 3982*delay_incr;
elsif nramp = '0' and StoredData = "111110001111" then SHout <= '1' after delay1 + 3983*delay_incr;
elsif nramp = '0' and StoredData = "111110010000" then SHout <= '1' after delay1 + 3984*delay_incr;
elsif nramp = '0' and StoredData = "111110010001" then SHout <= '1' after delay1 + 3985*delay_incr;
elsif nramp = '0' and StoredData = "111110010010" then SHout <= '1' after delay1 + 3986*delay_incr;
elsif nramp = '0' and StoredData = "111110010011" then SHout <= '1' after delay1 + 3987*delay_incr;
elsif nramp = '0' and StoredData = "111110010100" then SHout <= '1' after delay1 + 3988*delay_incr;
elsif nramp = '0' and StoredData = "111110010101" then SHout <= '1' after delay1 + 3989*delay_incr;
elsif nramp = '0' and StoredData = "111110010110" then SHout <= '1' after delay1 + 3990*delay_incr;
elsif nramp = '0' and StoredData = "111110010111" then SHout <= '1' after delay1 + 3991*delay_incr;
elsif nramp = '0' and StoredData = "111110011000" then SHout <= '1' after delay1 + 3992*delay_incr;
elsif nramp = '0' and StoredData = "111110011001" then SHout <= '1' after delay1 + 3993*delay_incr;
elsif nramp = '0' and StoredData = "111110011010" then SHout <= '1' after delay1 + 3994*delay_incr;
elsif nramp = '0' and StoredData = "111110011011" then SHout <= '1' after delay1 + 3995*delay_incr;
elsif nramp = '0' and StoredData = "111110011100" then SHout <= '1' after delay1 + 3996*delay_incr;
elsif nramp = '0' and StoredData = "111110011101" then SHout <= '1' after delay1 + 3997*delay_incr;
elsif nramp = '0' and StoredData = "111110011110" then SHout <= '1' after delay1 + 3998*delay_incr;
elsif nramp = '0' and StoredData = "111110011111" then SHout <= '1' after delay1 + 3999*delay_incr;
elsif nramp = '0' and StoredData = "111110100000" then SHout <= '1' after delay1 + 4000*delay_incr;
elsif nramp = '0' and StoredData = "111110100001" then SHout <= '1' after delay1 + 4001*delay_incr;
elsif nramp = '0' and StoredData = "111110100010" then SHout <= '1' after delay1 + 4002*delay_incr;
elsif nramp = '0' and StoredData = "111110100011" then SHout <= '1' after delay1 + 4003*delay_incr;
elsif nramp = '0' and StoredData = "111110100100" then SHout <= '1' after delay1 + 4004*delay_incr;
elsif nramp = '0' and StoredData = "111110100101" then SHout <= '1' after delay1 + 4005*delay_incr;
elsif nramp = '0' and StoredData = "111110100110" then SHout <= '1' after delay1 + 4006*delay_incr;
elsif nramp = '0' and StoredData = "111110100111" then SHout <= '1' after delay1 + 4007*delay_incr;
elsif nramp = '0' and StoredData = "111110101000" then SHout <= '1' after delay1 + 4008*delay_incr;
elsif nramp = '0' and StoredData = "111110101001" then SHout <= '1' after delay1 + 4009*delay_incr;
elsif nramp = '0' and StoredData = "111110101010" then SHout <= '1' after delay1 + 4010*delay_incr;
elsif nramp = '0' and StoredData = "111110101011" then SHout <= '1' after delay1 + 4011*delay_incr;
elsif nramp = '0' and StoredData = "111110101100" then SHout <= '1' after delay1 + 4012*delay_incr;
elsif nramp = '0' and StoredData = "111110101101" then SHout <= '1' after delay1 + 4013*delay_incr;
elsif nramp = '0' and StoredData = "111110101110" then SHout <= '1' after delay1 + 4014*delay_incr;
elsif nramp = '0' and StoredData = "111110101111" then SHout <= '1' after delay1 + 4015*delay_incr;
elsif nramp = '0' and StoredData = "111110110000" then SHout <= '1' after delay1 + 4016*delay_incr;
elsif nramp = '0' and StoredData = "111110110001" then SHout <= '1' after delay1 + 4017*delay_incr;
elsif nramp = '0' and StoredData = "111110110010" then SHout <= '1' after delay1 + 4018*delay_incr;
elsif nramp = '0' and StoredData = "111110110011" then SHout <= '1' after delay1 + 4019*delay_incr;
elsif nramp = '0' and StoredData = "111110110100" then SHout <= '1' after delay1 + 4020*delay_incr;
elsif nramp = '0' and StoredData = "111110110101" then SHout <= '1' after delay1 + 4021*delay_incr;
elsif nramp = '0' and StoredData = "111110110110" then SHout <= '1' after delay1 + 4022*delay_incr;
elsif nramp = '0' and StoredData = "111110110111" then SHout <= '1' after delay1 + 4023*delay_incr;
elsif nramp = '0' and StoredData = "111110111000" then SHout <= '1' after delay1 + 4024*delay_incr;
elsif nramp = '0' and StoredData = "111110111001" then SHout <= '1' after delay1 + 4025*delay_incr;
elsif nramp = '0' and StoredData = "111110111010" then SHout <= '1' after delay1 + 4026*delay_incr;
elsif nramp = '0' and StoredData = "111110111011" then SHout <= '1' after delay1 + 4027*delay_incr;
elsif nramp = '0' and StoredData = "111110111100" then SHout <= '1' after delay1 + 4028*delay_incr;
elsif nramp = '0' and StoredData = "111110111101" then SHout <= '1' after delay1 + 4029*delay_incr;
elsif nramp = '0' and StoredData = "111110111110" then SHout <= '1' after delay1 + 4030*delay_incr;
elsif nramp = '0' and StoredData = "111110111111" then SHout <= '1' after delay1 + 4031*delay_incr;
elsif nramp = '0' and StoredData = "111111000000" then SHout <= '1' after delay1 + 4032*delay_incr;
elsif nramp = '0' and StoredData = "111111000001" then SHout <= '1' after delay1 + 4033*delay_incr;
elsif nramp = '0' and StoredData = "111111000010" then SHout <= '1' after delay1 + 4034*delay_incr;
elsif nramp = '0' and StoredData = "111111000011" then SHout <= '1' after delay1 + 4035*delay_incr;
elsif nramp = '0' and StoredData = "111111000100" then SHout <= '1' after delay1 + 4036*delay_incr;
elsif nramp = '0' and StoredData = "111111000101" then SHout <= '1' after delay1 + 4037*delay_incr;
elsif nramp = '0' and StoredData = "111111000110" then SHout <= '1' after delay1 + 4038*delay_incr;
elsif nramp = '0' and StoredData = "111111000111" then SHout <= '1' after delay1 + 4039*delay_incr;
elsif nramp = '0' and StoredData = "111111001000" then SHout <= '1' after delay1 + 4040*delay_incr;
elsif nramp = '0' and StoredData = "111111001001" then SHout <= '1' after delay1 + 4041*delay_incr;
elsif nramp = '0' and StoredData = "111111001010" then SHout <= '1' after delay1 + 4042*delay_incr;
elsif nramp = '0' and StoredData = "111111001011" then SHout <= '1' after delay1 + 4043*delay_incr;
elsif nramp = '0' and StoredData = "111111001100" then SHout <= '1' after delay1 + 4044*delay_incr;
elsif nramp = '0' and StoredData = "111111001101" then SHout <= '1' after delay1 + 4045*delay_incr;
elsif nramp = '0' and StoredData = "111111001110" then SHout <= '1' after delay1 + 4046*delay_incr;
elsif nramp = '0' and StoredData = "111111001111" then SHout <= '1' after delay1 + 4047*delay_incr;
elsif nramp = '0' and StoredData = "111111010000" then SHout <= '1' after delay1 + 4048*delay_incr;
elsif nramp = '0' and StoredData = "111111010001" then SHout <= '1' after delay1 + 4049*delay_incr;
elsif nramp = '0' and StoredData = "111111010010" then SHout <= '1' after delay1 + 4050*delay_incr;
elsif nramp = '0' and StoredData = "111111010011" then SHout <= '1' after delay1 + 4051*delay_incr;
elsif nramp = '0' and StoredData = "111111010100" then SHout <= '1' after delay1 + 4052*delay_incr;
elsif nramp = '0' and StoredData = "111111010101" then SHout <= '1' after delay1 + 4053*delay_incr;
elsif nramp = '0' and StoredData = "111111010110" then SHout <= '1' after delay1 + 4054*delay_incr;
elsif nramp = '0' and StoredData = "111111010111" then SHout <= '1' after delay1 + 4055*delay_incr;
elsif nramp = '0' and StoredData = "111111011000" then SHout <= '1' after delay1 + 4056*delay_incr;
elsif nramp = '0' and StoredData = "111111011001" then SHout <= '1' after delay1 + 4057*delay_incr;
elsif nramp = '0' and StoredData = "111111011010" then SHout <= '1' after delay1 + 4058*delay_incr;
elsif nramp = '0' and StoredData = "111111011011" then SHout <= '1' after delay1 + 4059*delay_incr;
elsif nramp = '0' and StoredData = "111111011100" then SHout <= '1' after delay1 + 4060*delay_incr;
elsif nramp = '0' and StoredData = "111111011101" then SHout <= '1' after delay1 + 4061*delay_incr;
elsif nramp = '0' and StoredData = "111111011110" then SHout <= '1' after delay1 + 4062*delay_incr;
elsif nramp = '0' and StoredData = "111111011111" then SHout <= '1' after delay1 + 4063*delay_incr;
elsif nramp = '0' and StoredData = "111111100000" then SHout <= '1' after delay1 + 4064*delay_incr;
elsif nramp = '0' and StoredData = "111111100001" then SHout <= '1' after delay1 + 4065*delay_incr;
elsif nramp = '0' and StoredData = "111111100010" then SHout <= '1' after delay1 + 4066*delay_incr;
elsif nramp = '0' and StoredData = "111111100011" then SHout <= '1' after delay1 + 4067*delay_incr;
elsif nramp = '0' and StoredData = "111111100100" then SHout <= '1' after delay1 + 4068*delay_incr;
elsif nramp = '0' and StoredData = "111111100101" then SHout <= '1' after delay1 + 4069*delay_incr;
elsif nramp = '0' and StoredData = "111111100110" then SHout <= '1' after delay1 + 4070*delay_incr;
elsif nramp = '0' and StoredData = "111111100111" then SHout <= '1' after delay1 + 4071*delay_incr;
elsif nramp = '0' and StoredData = "111111101000" then SHout <= '1' after delay1 + 4072*delay_incr;
elsif nramp = '0' and StoredData = "111111101001" then SHout <= '1' after delay1 + 4073*delay_incr;
elsif nramp = '0' and StoredData = "111111101010" then SHout <= '1' after delay1 + 4074*delay_incr;
elsif nramp = '0' and StoredData = "111111101011" then SHout <= '1' after delay1 + 4075*delay_incr;
elsif nramp = '0' and StoredData = "111111101100" then SHout <= '1' after delay1 + 4076*delay_incr;
elsif nramp = '0' and StoredData = "111111101101" then SHout <= '1' after delay1 + 4077*delay_incr;
elsif nramp = '0' and StoredData = "111111101110" then SHout <= '1' after delay1 + 4078*delay_incr;
elsif nramp = '0' and StoredData = "111111101111" then SHout <= '1' after delay1 + 4079*delay_incr;
elsif nramp = '0' and StoredData = "111111110000" then SHout <= '1' after delay1 + 4080*delay_incr;
elsif nramp = '0' and StoredData = "111111110001" then SHout <= '1' after delay1 + 4081*delay_incr;
elsif nramp = '0' and StoredData = "111111110010" then SHout <= '1' after delay1 + 4082*delay_incr;
elsif nramp = '0' and StoredData = "111111110011" then SHout <= '1' after delay1 + 4083*delay_incr;
elsif nramp = '0' and StoredData = "111111110100" then SHout <= '1' after delay1 + 4084*delay_incr;
elsif nramp = '0' and StoredData = "111111110101" then SHout <= '1' after delay1 + 4085*delay_incr;
elsif nramp = '0' and StoredData = "111111110110" then SHout <= '1' after delay1 + 4086*delay_incr;
elsif nramp = '0' and StoredData = "111111110111" then SHout <= '1' after delay1 + 4087*delay_incr;
elsif nramp = '0' and StoredData = "111111111000" then SHout <= '1' after delay1 + 4088*delay_incr;
elsif nramp = '0' and StoredData = "111111111001" then SHout <= '1' after delay1 + 4089*delay_incr;
elsif nramp = '0' and StoredData = "111111111010" then SHout <= '1' after delay1 + 4090*delay_incr;
elsif nramp = '0' and StoredData = "111111111011" then SHout <= '1' after delay1 + 4091*delay_incr;
elsif nramp = '0' and StoredData = "111111111100" then SHout <= '1' after delay1 + 4092*delay_incr;
elsif nramp = '0' and StoredData = "111111111101" then SHout <= '1' after delay1 + 4093*delay_incr;
elsif nramp = '0' and StoredData = "111111111110" then SHout <= '1' after delay1 + 4094*delay_incr;
elsif nramp = '0' and StoredData = "111111111111" then SHout <= '1' after delay1 + 4095*delay_incr;
end if;
end process;
end behavioral;
